magic
tech sky130A
magscale 1 2
timestamp 1644002565
<< nwell >>
rect -48 3194 -30 3581
rect -48 2106 -32 2383
rect 504 697 520 1018
rect -48 -70 -30 180
rect -48 -1158 -32 -881
rect 504 -2567 520 -2246
rect -48 -3334 -30 -3084
rect -48 -4422 -32 -4145
rect 504 -5831 520 -5510
rect -48 -6598 -30 -6348
rect -48 -7686 -32 -7409
rect 504 -9095 520 -8774
rect -48 -9862 -30 -9612
rect -48 -10950 -32 -10673
rect 504 -12359 520 -12038
rect -48 -13126 -30 -12876
rect -48 -14214 -32 -13937
rect 504 -15623 520 -15302
rect -48 -16390 -30 -16140
rect -48 -17478 -32 -17201
rect 504 -18887 520 -18566
<< locali >>
rect 6262 963 6291 997
rect 6325 963 6383 997
rect 6417 963 6475 997
rect 6509 963 6567 997
rect 6601 963 6631 997
rect 541 581 575 701
rect 1504 651 1570 699
rect 6262 -2301 6291 -2267
rect 6325 -2301 6383 -2267
rect 6417 -2301 6475 -2267
rect 6509 -2301 6567 -2267
rect 6601 -2301 6631 -2267
rect 541 -2683 575 -2563
rect 1504 -2613 1570 -2565
rect 6262 -5565 6291 -5531
rect 6325 -5565 6383 -5531
rect 6417 -5565 6475 -5531
rect 6509 -5565 6567 -5531
rect 6601 -5565 6631 -5531
rect 541 -5947 575 -5827
rect 1504 -5877 1570 -5829
rect 6262 -8829 6291 -8795
rect 6325 -8829 6383 -8795
rect 6417 -8829 6475 -8795
rect 6509 -8829 6567 -8795
rect 6601 -8829 6631 -8795
rect 541 -9211 575 -9091
rect 1504 -9141 1570 -9093
rect 6262 -12093 6291 -12059
rect 6325 -12093 6383 -12059
rect 6417 -12093 6475 -12059
rect 6509 -12093 6567 -12059
rect 6601 -12093 6631 -12059
rect 541 -12475 575 -12355
rect 1504 -12405 1570 -12357
rect 6262 -15357 6291 -15323
rect 6325 -15357 6383 -15323
rect 6417 -15357 6475 -15323
rect 6509 -15357 6567 -15323
rect 6601 -15357 6631 -15323
rect 541 -15739 575 -15619
rect 1504 -15669 1570 -15621
rect 6262 -18621 6291 -18587
rect 6325 -18621 6383 -18587
rect 6417 -18621 6475 -18587
rect 6509 -18621 6567 -18587
rect 6601 -18621 6631 -18587
rect 541 -19003 575 -18883
rect 1504 -18933 1570 -18885
rect 6262 -19165 6291 -19131
rect 6325 -19165 6383 -19131
rect 6417 -19165 6475 -19131
rect 6509 -19165 6567 -19131
rect 6601 -19165 6631 -19131
<< viali >>
rect 262 3921 296 3955
rect 360 3921 394 3955
rect 538 3921 572 3955
rect 636 3921 670 3955
rect 813 3921 847 3955
rect 911 3921 945 3955
rect 1088 3921 1122 3955
rect 1186 3921 1220 3955
rect -431 3356 -395 3393
rect -249 2953 -198 3004
rect -249 2277 -198 2315
rect -245 1822 -204 1866
rect 6291 963 6325 997
rect 6383 963 6417 997
rect 6475 963 6509 997
rect 6567 963 6601 997
rect -145 656 -111 690
rect 24 656 58 690
rect -431 92 -395 129
rect -249 -311 -198 -260
rect -249 -987 -198 -949
rect -245 -1442 -204 -1398
rect 6291 -2301 6325 -2267
rect 6383 -2301 6417 -2267
rect 6475 -2301 6509 -2267
rect 6567 -2301 6601 -2267
rect -145 -2608 -111 -2574
rect 24 -2608 58 -2574
rect -431 -3172 -395 -3135
rect -249 -3575 -198 -3524
rect -249 -4251 -198 -4213
rect -245 -4706 -204 -4662
rect 6291 -5565 6325 -5531
rect 6383 -5565 6417 -5531
rect 6475 -5565 6509 -5531
rect 6567 -5565 6601 -5531
rect -145 -5872 -111 -5838
rect 24 -5872 58 -5838
rect -431 -6436 -395 -6399
rect -249 -6839 -198 -6788
rect -249 -7515 -198 -7477
rect -245 -7970 -204 -7926
rect 6291 -8829 6325 -8795
rect 6383 -8829 6417 -8795
rect 6475 -8829 6509 -8795
rect 6567 -8829 6601 -8795
rect -145 -9136 -111 -9102
rect 24 -9136 58 -9102
rect -431 -9700 -395 -9663
rect -249 -10103 -198 -10052
rect -249 -10779 -198 -10741
rect -245 -11234 -204 -11190
rect 6291 -12093 6325 -12059
rect 6383 -12093 6417 -12059
rect 6475 -12093 6509 -12059
rect 6567 -12093 6601 -12059
rect -145 -12400 -111 -12366
rect 24 -12400 58 -12366
rect -431 -12964 -395 -12927
rect -249 -13367 -198 -13316
rect -249 -14043 -198 -14005
rect -245 -14498 -204 -14454
rect 6291 -15357 6325 -15323
rect 6383 -15357 6417 -15323
rect 6475 -15357 6509 -15323
rect 6567 -15357 6601 -15323
rect -145 -15664 -111 -15630
rect 24 -15664 58 -15630
rect -431 -16228 -395 -16191
rect -249 -16631 -198 -16580
rect -249 -17307 -198 -17269
rect -245 -17762 -204 -17718
rect 6291 -18621 6325 -18587
rect 6383 -18621 6417 -18587
rect 6475 -18621 6509 -18587
rect 6567 -18621 6601 -18587
rect -145 -18928 -111 -18894
rect 24 -18928 58 -18894
rect 6291 -19165 6325 -19131
rect 6383 -19165 6417 -19131
rect 6475 -19165 6509 -19131
rect 6567 -19165 6601 -19131
<< metal1 >>
rect 6503 4222 6509 4280
rect 6567 4222 6573 4280
rect 240 3915 250 3980
rect 308 3915 318 3980
rect 346 3909 355 3980
rect 407 3909 417 3980
rect 516 3915 526 3980
rect 584 3915 594 3980
rect 622 3909 631 3980
rect 683 3909 692 3980
rect 791 3915 801 3980
rect 859 3915 869 3980
rect 897 3909 906 3980
rect 958 3909 967 3980
rect 1066 3915 1076 3980
rect 1134 3915 1144 3980
rect 1172 3909 1181 3980
rect 1233 3909 1242 3980
rect -437 3393 -389 3405
rect -437 3376 -431 3393
rect -395 3382 -389 3393
rect -395 3376 -385 3382
rect -437 3318 -385 3324
rect 345 3232 355 3284
rect 407 3232 417 3284
rect -248 3010 -181 3041
rect 621 3028 631 3080
rect 683 3028 693 3080
rect -261 3004 -181 3010
rect -261 2953 -249 3004
rect -198 2964 -181 3004
rect -261 2947 -248 2953
rect -248 2891 -181 2897
rect -400 2824 -394 2876
rect -342 2824 -336 2876
rect 896 2852 906 2904
rect 958 2852 968 2904
rect 1171 2772 1181 2824
rect 1233 2772 1243 2824
rect -400 2348 -394 2400
rect -342 2348 -336 2400
rect -254 2321 -248 2366
rect -261 2315 -248 2321
rect -181 2321 -175 2366
rect 78 2321 134 2385
rect -261 2277 -249 2315
rect -181 2299 134 2321
rect -198 2277 134 2299
rect -261 2271 134 2277
rect -251 1866 150 1878
rect -251 1822 -245 1866
rect -204 1822 150 1866
rect -251 1810 150 1822
rect -448 1731 -442 1793
rect -380 1731 -374 1793
rect 66 1781 150 1810
rect -432 1722 -389 1731
rect 1633 1390 1685 1396
rect 1743 1310 1753 1362
rect 1805 1310 1815 1362
rect 1863 1140 1873 1192
rect 1925 1140 1935 1192
rect 1983 1060 1993 1112
rect 2045 1060 2055 1112
rect 6262 1016 6631 1028
rect 6262 997 6509 1016
rect 6262 963 6291 997
rect 6325 963 6383 997
rect 6417 963 6475 997
rect 6262 958 6509 963
rect 6567 997 6631 1016
rect 6601 963 6631 997
rect 6567 958 6631 963
rect 6262 932 6631 958
rect -151 694 -105 696
rect 12 694 70 696
rect -165 690 70 694
rect -165 656 -145 690
rect -111 656 24 690
rect 58 656 70 690
rect -165 651 70 656
rect -151 650 -105 651
rect 12 650 70 651
rect -437 129 -389 141
rect -437 112 -431 129
rect -395 118 -389 129
rect -395 112 -385 118
rect -437 54 -385 60
rect 345 -32 355 20
rect 407 -32 417 20
rect -248 -254 -181 -223
rect 621 -236 631 -184
rect 683 -236 693 -184
rect -261 -260 -181 -254
rect -261 -311 -249 -260
rect -198 -300 -181 -260
rect -261 -317 -248 -311
rect -248 -373 -181 -367
rect -400 -440 -394 -388
rect -342 -440 -336 -388
rect 896 -412 906 -360
rect 958 -412 968 -360
rect 1171 -492 1181 -440
rect 1233 -492 1243 -440
rect -400 -916 -394 -864
rect -342 -916 -336 -864
rect -254 -943 -248 -898
rect -261 -949 -248 -943
rect -181 -943 -175 -898
rect 78 -943 134 -879
rect -261 -987 -249 -949
rect -181 -965 134 -943
rect -198 -987 134 -965
rect -261 -993 134 -987
rect -251 -1398 150 -1386
rect -251 -1442 -245 -1398
rect -204 -1442 150 -1398
rect -251 -1454 150 -1442
rect -448 -1533 -442 -1471
rect -380 -1533 -374 -1471
rect 66 -1483 150 -1454
rect -432 -1542 -389 -1533
rect 1623 -1874 1633 -1822
rect 1685 -1874 1695 -1822
rect 1743 -1954 1753 -1902
rect 1805 -1954 1815 -1902
rect 1863 -2124 1873 -2072
rect 1925 -2124 1935 -2072
rect 1983 -2204 1993 -2152
rect 2045 -2204 2055 -2152
rect 6262 -2248 6631 -2236
rect 6262 -2267 6509 -2248
rect 6262 -2301 6291 -2267
rect 6325 -2301 6383 -2267
rect 6417 -2301 6475 -2267
rect 6262 -2306 6509 -2301
rect 6567 -2267 6631 -2248
rect 6601 -2301 6631 -2267
rect 6567 -2306 6631 -2301
rect 6262 -2332 6631 -2306
rect -151 -2570 -105 -2568
rect 12 -2570 70 -2568
rect -165 -2574 70 -2570
rect -165 -2608 -145 -2574
rect -111 -2608 24 -2574
rect 58 -2608 70 -2574
rect -165 -2613 70 -2608
rect -151 -2614 -105 -2613
rect 12 -2614 70 -2613
rect -437 -3135 -389 -3123
rect -437 -3152 -431 -3135
rect -395 -3146 -389 -3135
rect -395 -3152 -385 -3146
rect -437 -3210 -385 -3204
rect 345 -3296 355 -3244
rect 407 -3296 417 -3244
rect -248 -3518 -181 -3487
rect 621 -3500 631 -3448
rect 683 -3500 693 -3448
rect -261 -3524 -181 -3518
rect -261 -3575 -249 -3524
rect -198 -3564 -181 -3524
rect -261 -3581 -248 -3575
rect -248 -3637 -181 -3631
rect -400 -3704 -394 -3652
rect -342 -3704 -336 -3652
rect 896 -3676 906 -3624
rect 958 -3676 968 -3624
rect 1171 -3756 1181 -3704
rect 1233 -3756 1243 -3704
rect -400 -4180 -394 -4128
rect -342 -4180 -336 -4128
rect -254 -4207 -248 -4162
rect -261 -4213 -248 -4207
rect -181 -4207 -175 -4162
rect 78 -4207 134 -4143
rect -261 -4251 -249 -4213
rect -181 -4229 134 -4207
rect -198 -4251 134 -4229
rect -261 -4257 134 -4251
rect -251 -4662 150 -4650
rect -251 -4706 -245 -4662
rect -204 -4706 150 -4662
rect -251 -4718 150 -4706
rect -448 -4797 -442 -4735
rect -380 -4797 -374 -4735
rect 66 -4747 150 -4718
rect -432 -4806 -389 -4797
rect 1623 -5132 1633 -5080
rect 1685 -5132 1695 -5080
rect 1743 -5218 1753 -5166
rect 1805 -5218 1815 -5166
rect 1863 -5388 1873 -5336
rect 1925 -5388 1935 -5336
rect 1983 -5468 1993 -5416
rect 2045 -5468 2055 -5416
rect 6262 -5512 6631 -5500
rect 6262 -5531 6509 -5512
rect 6262 -5565 6291 -5531
rect 6325 -5565 6383 -5531
rect 6417 -5565 6475 -5531
rect 6262 -5570 6509 -5565
rect 6567 -5531 6631 -5512
rect 6601 -5565 6631 -5531
rect 6567 -5570 6631 -5565
rect 6262 -5596 6631 -5570
rect -151 -5834 -105 -5832
rect 12 -5834 70 -5832
rect -165 -5838 70 -5834
rect -165 -5872 -145 -5838
rect -111 -5872 24 -5838
rect 58 -5872 70 -5838
rect -165 -5877 70 -5872
rect -151 -5878 -105 -5877
rect 12 -5878 70 -5877
rect -437 -6399 -389 -6387
rect -437 -6416 -431 -6399
rect -395 -6410 -389 -6399
rect -395 -6416 -385 -6410
rect -437 -6474 -385 -6468
rect 345 -6560 355 -6508
rect 407 -6560 417 -6508
rect -248 -6782 -181 -6751
rect 621 -6764 631 -6712
rect 683 -6764 693 -6712
rect -261 -6788 -181 -6782
rect -261 -6839 -249 -6788
rect -198 -6828 -181 -6788
rect -261 -6845 -248 -6839
rect -248 -6901 -181 -6895
rect -400 -6968 -394 -6916
rect -342 -6968 -336 -6916
rect 896 -6940 906 -6888
rect 958 -6940 968 -6888
rect 1171 -7020 1181 -6968
rect 1233 -7020 1243 -6968
rect -400 -7444 -394 -7392
rect -342 -7444 -336 -7392
rect -254 -7471 -248 -7426
rect -261 -7477 -248 -7471
rect -181 -7471 -175 -7426
rect 78 -7471 134 -7407
rect -261 -7515 -249 -7477
rect -181 -7493 134 -7471
rect -198 -7515 134 -7493
rect -261 -7521 134 -7515
rect -251 -7926 150 -7914
rect -251 -7970 -245 -7926
rect -204 -7970 150 -7926
rect -251 -7982 150 -7970
rect -448 -8061 -442 -7999
rect -380 -8061 -374 -7999
rect 66 -8011 150 -7982
rect -432 -8070 -389 -8061
rect 1623 -8396 1633 -8344
rect 1685 -8396 1695 -8344
rect 1743 -8482 1753 -8430
rect 1805 -8482 1815 -8430
rect 1863 -8652 1873 -8600
rect 1925 -8652 1935 -8600
rect 1983 -8732 1993 -8680
rect 2045 -8732 2055 -8680
rect 6262 -8776 6631 -8764
rect 6262 -8795 6509 -8776
rect 6262 -8829 6291 -8795
rect 6325 -8829 6383 -8795
rect 6417 -8829 6475 -8795
rect 6262 -8834 6509 -8829
rect 6567 -8795 6631 -8776
rect 6601 -8829 6631 -8795
rect 6567 -8834 6631 -8829
rect 6262 -8860 6631 -8834
rect -151 -9098 -105 -9096
rect 12 -9098 70 -9096
rect -165 -9102 70 -9098
rect -165 -9136 -145 -9102
rect -111 -9136 24 -9102
rect 58 -9136 70 -9102
rect -165 -9141 70 -9136
rect -151 -9142 -105 -9141
rect 12 -9142 70 -9141
rect -437 -9663 -389 -9651
rect -437 -9680 -431 -9663
rect -395 -9674 -389 -9663
rect -395 -9680 -385 -9674
rect -437 -9738 -385 -9732
rect 345 -9824 355 -9772
rect 407 -9824 417 -9772
rect -248 -10046 -181 -10015
rect 621 -10028 631 -9976
rect 683 -10028 693 -9976
rect -261 -10052 -181 -10046
rect -261 -10103 -249 -10052
rect -198 -10092 -181 -10052
rect -261 -10109 -248 -10103
rect -248 -10165 -181 -10159
rect -400 -10232 -394 -10180
rect -342 -10232 -336 -10180
rect 896 -10204 906 -10152
rect 958 -10204 968 -10152
rect 1171 -10284 1181 -10232
rect 1233 -10284 1243 -10232
rect -400 -10708 -394 -10656
rect -342 -10708 -336 -10656
rect -254 -10735 -248 -10690
rect -261 -10741 -248 -10735
rect -181 -10735 -175 -10690
rect 78 -10735 134 -10671
rect -261 -10779 -249 -10741
rect -181 -10757 134 -10735
rect -198 -10779 134 -10757
rect -261 -10785 134 -10779
rect -251 -11190 150 -11178
rect -251 -11234 -245 -11190
rect -204 -11234 150 -11190
rect -251 -11246 150 -11234
rect -448 -11325 -442 -11263
rect -380 -11325 -374 -11263
rect 66 -11275 150 -11246
rect -432 -11334 -389 -11325
rect 1623 -11660 1633 -11608
rect 1685 -11660 1695 -11608
rect 1743 -11746 1753 -11694
rect 1805 -11746 1815 -11694
rect 1863 -11916 1873 -11864
rect 1925 -11916 1935 -11864
rect 1983 -11996 1993 -11944
rect 2045 -11996 2055 -11944
rect 6262 -12040 6631 -12028
rect 6262 -12059 6509 -12040
rect 6262 -12093 6291 -12059
rect 6325 -12093 6383 -12059
rect 6417 -12093 6475 -12059
rect 6262 -12098 6509 -12093
rect 6567 -12059 6631 -12040
rect 6601 -12093 6631 -12059
rect 6567 -12098 6631 -12093
rect 6262 -12124 6631 -12098
rect -151 -12362 -105 -12360
rect 12 -12362 70 -12360
rect -165 -12366 70 -12362
rect -165 -12400 -145 -12366
rect -111 -12400 24 -12366
rect 58 -12400 70 -12366
rect -165 -12405 70 -12400
rect -151 -12406 -105 -12405
rect 12 -12406 70 -12405
rect -437 -12927 -389 -12915
rect -437 -12944 -431 -12927
rect -395 -12938 -389 -12927
rect -395 -12944 -385 -12938
rect -437 -13002 -385 -12996
rect 345 -13088 355 -13036
rect 407 -13088 417 -13036
rect -248 -13310 -181 -13279
rect 621 -13292 631 -13240
rect 683 -13292 693 -13240
rect -261 -13316 -181 -13310
rect -261 -13367 -249 -13316
rect -198 -13356 -181 -13316
rect -261 -13373 -248 -13367
rect -248 -13429 -181 -13423
rect -400 -13496 -394 -13444
rect -342 -13496 -336 -13444
rect 896 -13468 906 -13416
rect 958 -13468 968 -13416
rect 1171 -13548 1181 -13496
rect 1233 -13548 1243 -13496
rect -400 -13972 -394 -13920
rect -342 -13972 -336 -13920
rect -254 -13999 -248 -13954
rect -261 -14005 -248 -13999
rect -181 -13999 -175 -13954
rect 78 -13999 134 -13935
rect -261 -14043 -249 -14005
rect -181 -14021 134 -13999
rect -198 -14043 134 -14021
rect -261 -14049 134 -14043
rect -251 -14454 150 -14442
rect -251 -14498 -245 -14454
rect -204 -14498 150 -14454
rect -251 -14510 150 -14498
rect -448 -14589 -442 -14527
rect -380 -14589 -374 -14527
rect 66 -14539 150 -14510
rect -432 -14598 -389 -14589
rect 1623 -14924 1633 -14872
rect 1685 -14924 1695 -14872
rect 1743 -15010 1753 -14958
rect 1805 -15010 1815 -14958
rect 1863 -15180 1873 -15128
rect 1925 -15180 1935 -15128
rect 1983 -15260 1993 -15208
rect 2045 -15260 2055 -15208
rect 6262 -15304 6631 -15292
rect 6262 -15323 6509 -15304
rect 6262 -15357 6291 -15323
rect 6325 -15357 6383 -15323
rect 6417 -15357 6475 -15323
rect 6262 -15362 6509 -15357
rect 6567 -15323 6631 -15304
rect 6601 -15357 6631 -15323
rect 6567 -15362 6631 -15357
rect 6262 -15388 6631 -15362
rect -151 -15626 -105 -15624
rect 12 -15626 70 -15624
rect -165 -15630 70 -15626
rect -165 -15664 -145 -15630
rect -111 -15664 24 -15630
rect 58 -15664 70 -15630
rect -165 -15669 70 -15664
rect -151 -15670 -105 -15669
rect 12 -15670 70 -15669
rect -437 -16191 -389 -16179
rect -437 -16208 -431 -16191
rect -395 -16202 -389 -16191
rect -395 -16208 -385 -16202
rect -437 -16266 -385 -16260
rect 345 -16352 355 -16300
rect 407 -16352 417 -16300
rect -248 -16574 -181 -16543
rect 621 -16556 631 -16504
rect 683 -16556 693 -16504
rect -261 -16580 -181 -16574
rect -261 -16631 -249 -16580
rect -198 -16620 -181 -16580
rect -261 -16637 -248 -16631
rect -248 -16693 -181 -16687
rect -400 -16760 -394 -16708
rect -342 -16760 -336 -16708
rect 896 -16732 906 -16680
rect 958 -16732 968 -16680
rect 1171 -16812 1181 -16760
rect 1233 -16812 1243 -16760
rect -400 -17236 -394 -17184
rect -342 -17236 -336 -17184
rect -254 -17263 -248 -17218
rect -261 -17269 -248 -17263
rect -181 -17263 -175 -17218
rect 78 -17263 134 -17199
rect -261 -17307 -249 -17269
rect -181 -17285 134 -17263
rect -198 -17307 134 -17285
rect -261 -17313 134 -17307
rect -251 -17718 150 -17706
rect -251 -17762 -245 -17718
rect -204 -17762 150 -17718
rect -251 -17774 150 -17762
rect -448 -17853 -442 -17791
rect -380 -17853 -374 -17791
rect 66 -17803 150 -17774
rect -432 -17862 -389 -17853
rect 1623 -18188 1633 -18136
rect 1685 -18188 1695 -18136
rect 1743 -18274 1753 -18222
rect 1805 -18274 1815 -18222
rect 1863 -18444 1873 -18392
rect 1925 -18444 1935 -18392
rect 1983 -18524 1993 -18472
rect 2045 -18524 2055 -18472
rect 6262 -18568 6631 -18556
rect 6262 -18587 6509 -18568
rect 6262 -18621 6291 -18587
rect 6325 -18621 6383 -18587
rect 6417 -18621 6475 -18587
rect 6262 -18626 6509 -18621
rect 6567 -18587 6631 -18568
rect 6601 -18621 6631 -18587
rect 6567 -18626 6631 -18621
rect 6262 -18652 6631 -18626
rect -151 -18890 -105 -18888
rect 12 -18890 70 -18888
rect -165 -18894 70 -18890
rect -165 -18928 -145 -18894
rect -111 -18928 24 -18894
rect 58 -18928 70 -18894
rect -165 -18933 70 -18928
rect -151 -18934 -105 -18933
rect 12 -18934 70 -18933
rect 6262 -19112 6631 -19100
rect 6262 -19131 6409 -19112
rect 6467 -19131 6631 -19112
rect 6262 -19165 6291 -19131
rect 6325 -19165 6383 -19131
rect 6467 -19165 6475 -19131
rect 6509 -19165 6567 -19131
rect 6601 -19165 6631 -19131
rect 6262 -19170 6409 -19165
rect 6467 -19170 6631 -19165
rect 6262 -19196 6631 -19170
<< via1 >>
rect 6509 4222 6567 4280
rect 250 3955 308 3980
rect 250 3921 262 3955
rect 262 3921 296 3955
rect 296 3921 308 3955
rect 250 3915 308 3921
rect 355 3955 407 3980
rect 355 3921 360 3955
rect 360 3921 394 3955
rect 394 3921 407 3955
rect 355 3909 407 3921
rect 526 3955 584 3980
rect 526 3921 538 3955
rect 538 3921 572 3955
rect 572 3921 584 3955
rect 526 3915 584 3921
rect 631 3955 683 3980
rect 631 3921 636 3955
rect 636 3921 670 3955
rect 670 3921 683 3955
rect 631 3909 683 3921
rect 801 3955 859 3980
rect 801 3921 813 3955
rect 813 3921 847 3955
rect 847 3921 859 3955
rect 801 3915 859 3921
rect 906 3955 958 3980
rect 906 3921 911 3955
rect 911 3921 945 3955
rect 945 3921 958 3955
rect 906 3909 958 3921
rect 1076 3955 1134 3980
rect 1076 3921 1088 3955
rect 1088 3921 1122 3955
rect 1122 3921 1134 3955
rect 1076 3915 1134 3921
rect 1181 3955 1233 3980
rect 1181 3921 1186 3955
rect 1186 3921 1220 3955
rect 1220 3921 1233 3955
rect 1181 3909 1233 3921
rect 6409 3678 6467 3736
rect -437 3356 -431 3376
rect -431 3356 -395 3376
rect -395 3356 -385 3376
rect -437 3324 -385 3356
rect 355 3232 407 3284
rect 6509 3134 6567 3192
rect 631 3028 683 3080
rect -248 2953 -198 2964
rect -198 2953 -181 2964
rect -248 2897 -181 2953
rect -394 2824 -342 2876
rect 906 2852 958 2904
rect 1181 2772 1233 2824
rect 6409 2590 6467 2648
rect -394 2348 -342 2400
rect -248 2315 -181 2366
rect -248 2299 -198 2315
rect -198 2299 -181 2315
rect 6509 2046 6567 2104
rect -442 1731 -380 1793
rect 6409 1502 6467 1560
rect 1633 1396 1685 1448
rect 1753 1310 1805 1362
rect 1873 1140 1925 1192
rect 1993 1060 2045 1112
rect 6509 958 6567 1016
rect 6409 414 6467 472
rect -437 92 -431 112
rect -431 92 -395 112
rect -395 92 -385 112
rect -437 60 -385 92
rect 355 -32 407 20
rect 6509 -130 6567 -72
rect 631 -236 683 -184
rect -248 -311 -198 -300
rect -198 -311 -181 -300
rect -248 -367 -181 -311
rect -394 -440 -342 -388
rect 906 -412 958 -360
rect 1181 -492 1233 -440
rect 6409 -674 6467 -616
rect -394 -916 -342 -864
rect -248 -949 -181 -898
rect -248 -965 -198 -949
rect -198 -965 -181 -949
rect 6509 -1218 6567 -1160
rect -442 -1533 -380 -1471
rect 6409 -1762 6467 -1704
rect 1633 -1874 1685 -1822
rect 1753 -1954 1805 -1902
rect 1873 -2124 1925 -2072
rect 1993 -2204 2045 -2152
rect 6509 -2306 6567 -2248
rect 6409 -2850 6467 -2792
rect -437 -3172 -431 -3152
rect -431 -3172 -395 -3152
rect -395 -3172 -385 -3152
rect -437 -3204 -385 -3172
rect 355 -3296 407 -3244
rect 6509 -3394 6567 -3336
rect 631 -3500 683 -3448
rect -248 -3575 -198 -3564
rect -198 -3575 -181 -3564
rect -248 -3631 -181 -3575
rect -394 -3704 -342 -3652
rect 906 -3676 958 -3624
rect 1181 -3756 1233 -3704
rect 6409 -3938 6467 -3880
rect -394 -4180 -342 -4128
rect -248 -4213 -181 -4162
rect -248 -4229 -198 -4213
rect -198 -4229 -181 -4213
rect 6509 -4482 6567 -4424
rect -442 -4797 -380 -4735
rect 6409 -5026 6467 -4968
rect 1633 -5132 1685 -5080
rect 1753 -5218 1805 -5166
rect 1873 -5388 1925 -5336
rect 1993 -5468 2045 -5416
rect 6509 -5570 6567 -5512
rect 6409 -6114 6467 -6056
rect -437 -6436 -431 -6416
rect -431 -6436 -395 -6416
rect -395 -6436 -385 -6416
rect -437 -6468 -385 -6436
rect 355 -6560 407 -6508
rect 6509 -6658 6567 -6600
rect 631 -6764 683 -6712
rect -248 -6839 -198 -6828
rect -198 -6839 -181 -6828
rect -248 -6895 -181 -6839
rect -394 -6968 -342 -6916
rect 906 -6940 958 -6888
rect 1181 -7020 1233 -6968
rect 6409 -7202 6467 -7144
rect -394 -7444 -342 -7392
rect -248 -7477 -181 -7426
rect -248 -7493 -198 -7477
rect -198 -7493 -181 -7477
rect 6509 -7746 6567 -7688
rect -442 -8061 -380 -7999
rect 6409 -8290 6467 -8232
rect 1633 -8396 1685 -8344
rect 1753 -8482 1805 -8430
rect 1873 -8652 1925 -8600
rect 1993 -8732 2045 -8680
rect 6509 -8834 6567 -8776
rect 6409 -9378 6467 -9320
rect -437 -9700 -431 -9680
rect -431 -9700 -395 -9680
rect -395 -9700 -385 -9680
rect -437 -9732 -385 -9700
rect 355 -9824 407 -9772
rect 6509 -9922 6567 -9864
rect 631 -10028 683 -9976
rect -248 -10103 -198 -10092
rect -198 -10103 -181 -10092
rect -248 -10159 -181 -10103
rect -394 -10232 -342 -10180
rect 906 -10204 958 -10152
rect 1181 -10284 1233 -10232
rect 6409 -10466 6467 -10408
rect -394 -10708 -342 -10656
rect -248 -10741 -181 -10690
rect -248 -10757 -198 -10741
rect -198 -10757 -181 -10741
rect 6509 -11010 6567 -10952
rect -442 -11325 -380 -11263
rect 6409 -11554 6467 -11496
rect 1633 -11660 1685 -11608
rect 1753 -11746 1805 -11694
rect 1873 -11916 1925 -11864
rect 1993 -11996 2045 -11944
rect 6509 -12098 6567 -12040
rect 6409 -12642 6467 -12584
rect -437 -12964 -431 -12944
rect -431 -12964 -395 -12944
rect -395 -12964 -385 -12944
rect -437 -12996 -385 -12964
rect 355 -13088 407 -13036
rect 6509 -13186 6567 -13128
rect 631 -13292 683 -13240
rect -248 -13367 -198 -13356
rect -198 -13367 -181 -13356
rect -248 -13423 -181 -13367
rect -394 -13496 -342 -13444
rect 906 -13468 958 -13416
rect 1181 -13548 1233 -13496
rect 6409 -13730 6467 -13672
rect -394 -13972 -342 -13920
rect -248 -14005 -181 -13954
rect -248 -14021 -198 -14005
rect -198 -14021 -181 -14005
rect 6509 -14274 6567 -14216
rect -442 -14589 -380 -14527
rect 6409 -14818 6467 -14760
rect 1633 -14924 1685 -14872
rect 1753 -15010 1805 -14958
rect 1873 -15180 1925 -15128
rect 1993 -15260 2045 -15208
rect 6509 -15362 6567 -15304
rect 6409 -15906 6467 -15848
rect -437 -16228 -431 -16208
rect -431 -16228 -395 -16208
rect -395 -16228 -385 -16208
rect -437 -16260 -385 -16228
rect 355 -16352 407 -16300
rect 6509 -16450 6567 -16392
rect 631 -16556 683 -16504
rect -248 -16631 -198 -16620
rect -198 -16631 -181 -16620
rect -248 -16687 -181 -16631
rect -394 -16760 -342 -16708
rect 906 -16732 958 -16680
rect 1181 -16812 1233 -16760
rect 6409 -16994 6467 -16936
rect -394 -17236 -342 -17184
rect -248 -17269 -181 -17218
rect -248 -17285 -198 -17269
rect -198 -17285 -181 -17269
rect 6509 -17538 6567 -17480
rect -442 -17853 -380 -17791
rect 6409 -18082 6467 -18024
rect 1633 -18188 1685 -18136
rect 1753 -18274 1805 -18222
rect 1873 -18444 1925 -18392
rect 1993 -18524 2045 -18472
rect 6509 -18626 6567 -18568
rect 6409 -19131 6467 -19112
rect 6409 -19165 6417 -19131
rect 6417 -19165 6467 -19131
rect 6409 -19170 6467 -19165
<< metal2 >>
rect 250 3980 308 4292
rect 250 3905 308 3915
rect 355 3980 407 3990
rect -442 3376 -380 3381
rect -443 3324 -437 3376
rect -385 3324 -379 3376
rect -442 2882 -380 3324
rect 355 3284 407 3909
rect 526 3980 584 4292
rect 526 3905 584 3915
rect 631 3980 683 3990
rect -254 2897 -248 2964
rect -181 2897 -175 2964
rect -442 2876 -342 2882
rect -442 2824 -394 2876
rect -442 2818 -342 2824
rect -442 2406 -380 2818
rect -442 2400 -342 2406
rect -442 2348 -394 2400
rect -442 2342 -342 2348
rect -248 2366 -181 2897
rect -442 1793 -380 2342
rect -248 2265 -181 2299
rect -442 1725 -380 1731
rect -442 112 -380 117
rect -443 60 -437 112
rect -385 60 -379 112
rect -442 -382 -380 60
rect 355 20 407 3232
rect -254 -367 -248 -300
rect -181 -367 -175 -300
rect -442 -388 -342 -382
rect -442 -440 -394 -388
rect -442 -446 -342 -440
rect -442 -858 -380 -446
rect -442 -864 -342 -858
rect -442 -916 -394 -864
rect -442 -922 -342 -916
rect -248 -898 -181 -367
rect -442 -1471 -380 -922
rect -248 -999 -181 -965
rect -442 -1539 -380 -1533
rect -442 -3152 -380 -3147
rect -443 -3204 -437 -3152
rect -385 -3204 -379 -3152
rect -442 -3646 -380 -3204
rect 355 -3244 407 -32
rect -254 -3631 -248 -3564
rect -181 -3631 -175 -3564
rect -442 -3652 -342 -3646
rect -442 -3704 -394 -3652
rect -442 -3710 -342 -3704
rect -442 -4122 -380 -3710
rect -442 -4128 -342 -4122
rect -442 -4180 -394 -4128
rect -442 -4186 -342 -4180
rect -248 -4162 -181 -3631
rect -442 -4735 -380 -4186
rect -248 -4263 -181 -4229
rect -442 -4803 -380 -4797
rect -442 -6416 -380 -6411
rect -443 -6468 -437 -6416
rect -385 -6468 -379 -6416
rect -442 -6910 -380 -6468
rect 355 -6508 407 -3296
rect -254 -6895 -248 -6828
rect -181 -6895 -175 -6828
rect -442 -6916 -342 -6910
rect -442 -6968 -394 -6916
rect -442 -6974 -342 -6968
rect -442 -7386 -380 -6974
rect -442 -7392 -342 -7386
rect -442 -7444 -394 -7392
rect -442 -7450 -342 -7444
rect -248 -7426 -181 -6895
rect -442 -7999 -380 -7450
rect -248 -7527 -181 -7493
rect -442 -8067 -380 -8061
rect -442 -9680 -380 -9675
rect -443 -9732 -437 -9680
rect -385 -9732 -379 -9680
rect -442 -10174 -380 -9732
rect 355 -9772 407 -6560
rect -254 -10159 -248 -10092
rect -181 -10159 -175 -10092
rect -442 -10180 -342 -10174
rect -442 -10232 -394 -10180
rect -442 -10238 -342 -10232
rect -442 -10650 -380 -10238
rect -442 -10656 -342 -10650
rect -442 -10708 -394 -10656
rect -442 -10714 -342 -10708
rect -248 -10690 -181 -10159
rect -442 -11263 -380 -10714
rect -248 -10791 -181 -10757
rect -442 -11331 -380 -11325
rect -442 -12944 -380 -12939
rect -443 -12996 -437 -12944
rect -385 -12996 -379 -12944
rect -442 -13438 -380 -12996
rect 355 -13036 407 -9824
rect -254 -13423 -248 -13356
rect -181 -13423 -175 -13356
rect -442 -13444 -342 -13438
rect -442 -13496 -394 -13444
rect -442 -13502 -342 -13496
rect -442 -13914 -380 -13502
rect -442 -13920 -342 -13914
rect -442 -13972 -394 -13920
rect -442 -13978 -342 -13972
rect -248 -13954 -181 -13423
rect -442 -14527 -380 -13978
rect -248 -14055 -181 -14021
rect -442 -14595 -380 -14589
rect -442 -16208 -380 -16203
rect -443 -16260 -437 -16208
rect -385 -16260 -379 -16208
rect -442 -16702 -380 -16260
rect 355 -16300 407 -13088
rect 355 -16362 407 -16352
rect 631 3080 683 3909
rect 801 3980 859 4292
rect 801 3905 859 3915
rect 906 3980 958 3990
rect 631 -184 683 3028
rect 631 -3448 683 -236
rect 631 -6712 683 -3500
rect 631 -9976 683 -6764
rect 631 -13240 683 -10028
rect 631 -16504 683 -13292
rect 631 -16562 683 -16556
rect 906 2904 958 3909
rect 1076 3980 1134 4292
rect 1076 3905 1134 3915
rect 1181 3980 1233 3990
rect 906 -360 958 2852
rect 906 -3624 958 -412
rect 906 -6888 958 -3676
rect 906 -10152 958 -6940
rect 906 -13416 958 -10204
rect -254 -16687 -248 -16620
rect -181 -16687 -175 -16620
rect 906 -16680 958 -13468
rect -442 -16708 -342 -16702
rect -442 -16760 -394 -16708
rect -442 -16766 -342 -16760
rect -442 -17178 -380 -16766
rect -442 -17184 -342 -17178
rect -442 -17236 -394 -17184
rect -442 -17242 -342 -17236
rect -248 -17218 -181 -16687
rect 906 -16747 958 -16732
rect 1181 2824 1233 3909
rect 1181 -440 1233 2772
rect 1181 -3704 1233 -492
rect 1181 -6968 1233 -3756
rect 1181 -10232 1233 -7020
rect 1181 -13496 1233 -10284
rect 1181 -16760 1233 -13548
rect 1181 -16822 1233 -16812
rect 1633 3980 1691 4292
rect 1753 3980 1811 4292
rect 1873 3980 1931 4292
rect 1993 3980 2051 4292
rect 6509 4280 6567 4286
rect 1633 1448 1685 3980
rect 1633 -1822 1685 1396
rect 1633 -5080 1685 -1874
rect 1633 -8344 1685 -5132
rect 1633 -11608 1685 -8396
rect 1633 -14872 1685 -11660
rect -442 -17791 -380 -17242
rect -248 -17319 -181 -17285
rect -442 -17859 -380 -17853
rect 1633 -18136 1685 -14924
rect 1633 -18610 1685 -18188
rect 1753 1362 1805 3980
rect 1753 -1902 1805 1310
rect 1753 -5166 1805 -1954
rect 1753 -8430 1805 -5218
rect 1753 -11694 1805 -8482
rect 1753 -14958 1805 -11746
rect 1753 -18222 1805 -15010
rect 1753 -18610 1805 -18274
rect 1873 1192 1925 3980
rect 1873 -2072 1925 1140
rect 1873 -5336 1925 -2124
rect 1873 -8600 1925 -5388
rect 1873 -11864 1925 -8652
rect 1873 -15128 1925 -11916
rect 1873 -18392 1925 -15180
rect 1873 -18610 1925 -18444
rect 1993 1112 2045 3980
rect 6409 3736 6467 3742
rect 1993 -2152 2045 1060
rect 1993 -5416 2045 -2204
rect 1993 -8680 2045 -5468
rect 1993 -11944 2045 -8732
rect 1993 -15208 2045 -11996
rect 1993 -18472 2045 -15260
rect 1993 -18610 2045 -18524
rect 3696 -18799 3785 3396
rect 6409 2648 6467 3678
rect 6409 1560 6467 2590
rect 6409 472 6467 1502
rect 6409 -616 6467 414
rect 6409 -1704 6467 -674
rect 6409 -2792 6467 -1762
rect 6409 -3880 6467 -2850
rect 6409 -4968 6467 -3938
rect 6409 -6056 6467 -5026
rect 6409 -7144 6467 -6114
rect 6409 -8232 6467 -7202
rect 6409 -9320 6467 -8290
rect 6409 -10408 6467 -9378
rect 6409 -11496 6467 -10466
rect 6409 -12584 6467 -11554
rect 6409 -13672 6467 -12642
rect 6409 -14760 6467 -13730
rect 6409 -15848 6467 -14818
rect 6409 -16936 6467 -15906
rect 6409 -18024 6467 -16994
rect 6409 -19112 6467 -18082
rect 6509 3192 6567 4222
rect 6509 2104 6567 3134
rect 6509 1016 6567 2046
rect 6509 -72 6567 958
rect 6509 -1160 6567 -130
rect 6509 -2248 6567 -1218
rect 6509 -3336 6567 -2306
rect 6509 -4424 6567 -3394
rect 6509 -5512 6567 -4482
rect 6509 -6600 6567 -5570
rect 6509 -7688 6567 -6658
rect 6509 -8776 6567 -7746
rect 6509 -9864 6567 -8834
rect 6509 -10952 6567 -9922
rect 6509 -12040 6567 -11010
rect 6509 -13128 6567 -12098
rect 6509 -14216 6567 -13186
rect 6509 -15304 6567 -14274
rect 6509 -16392 6567 -15362
rect 6509 -17480 6567 -16450
rect 6509 -18568 6567 -17538
rect 6509 -18632 6567 -18626
rect 6409 -19176 6467 -19170
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_21 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1633901636
transform 1 0 -86 0 1 -18060
box -38 -48 130 592
use sky130_fd_sc_hd__clkinv_16  sky130_fd_sc_hd__clkinv_16_18 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1633901636
transform 1 0 -2294 0 1 -18060
box -38 -48 2246 592
use sky130_fd_sc_hd__clkinv_4  sky130_fd_sc_hd__clkinv_4_12 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1633901636
transform 1 0 -86 0 1 -19148
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_4  sky130_fd_sc_hd__clkinv_4_13
timestamp 1633901636
transform 1 0 -730 0 1 -19148
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_7
timestamp 1633901636
transform 1 0 -2294 0 1 -19148
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_8  sky130_fd_sc_hd__clkbuf_8_6 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1633901636
transform 1 0 558 0 1 -19148
box -38 -48 1050 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1633901636
transform 1 0 -2202 0 1 -19148
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_26
timestamp 1633901636
transform 1 0 -1466 0 1 -19148
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_20
timestamp 1633901636
transform 1 0 -86 0 1 -16972
box -38 -48 130 592
use sky130_fd_sc_hd__clkinv_16  sky130_fd_sc_hd__clkinv_16_19
timestamp 1633901636
transform 1 0 -2294 0 -1 -16972
box -38 -48 2246 592
use sky130_fd_sc_hd__clkinv_16  sky130_fd_sc_hd__clkinv_16_20
timestamp 1633901636
transform 1 0 -2294 0 1 -16972
box -38 -48 2246 592
use n-leg  n-leg_6
timestamp 1643392248
transform 1 0 -284 0 1 -19148
box 1854 -48 6546 1136
use p-leg  p-leg_6
timestamp 1643671812
transform 1 0 2 0 1 -18070
box -34 -38 6666 2234
use sky130_fd_sc_hd__clkinv_4  sky130_fd_sc_hd__clkinv_4_10
timestamp 1633901636
transform 1 0 -86 0 1 -15884
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_4  sky130_fd_sc_hd__clkinv_4_11
timestamp 1633901636
transform 1 0 -730 0 1 -15884
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_6
timestamp 1633901636
transform 1 0 -2294 0 1 -15884
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_16  sky130_fd_sc_hd__clkbuf_16_6 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1633901636
transform 1 0 -1926 0 -1 -15884
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_8  sky130_fd_sc_hd__clkbuf_8_5
timestamp 1633901636
transform 1 0 558 0 1 -15884
box -38 -48 1050 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_25
timestamp 1633901636
transform 1 0 -2202 0 1 -15884
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_24
timestamp 1633901636
transform 1 0 -1466 0 1 -15884
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_19
timestamp 1633901636
transform 1 0 -86 0 1 -14796
box -38 -48 130 592
use sky130_fd_sc_hd__clkinv_16  sky130_fd_sc_hd__clkinv_16_15
timestamp 1633901636
transform 1 0 -2294 0 1 -14796
box -38 -48 2246 592
use n-leg  n-leg_5
timestamp 1643392248
transform 1 0 -284 0 1 -15884
box 1854 -48 6546 1136
use p-leg  p-leg_5
timestamp 1643671812
transform 1 0 2 0 1 -14806
box -34 -38 6666 2234
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_18
timestamp 1633901636
transform 1 0 -86 0 1 -13708
box -38 -48 130 592
use sky130_fd_sc_hd__clkinv_16  sky130_fd_sc_hd__clkinv_16_17
timestamp 1633901636
transform 1 0 -2294 0 1 -13708
box -38 -48 2246 592
use sky130_fd_sc_hd__clkinv_16  sky130_fd_sc_hd__clkinv_16_16
timestamp 1633901636
transform 1 0 -2294 0 -1 -13708
box -38 -48 2246 592
use sky130_fd_sc_hd__clkinv_4  sky130_fd_sc_hd__clkinv_4_8
timestamp 1633901636
transform 1 0 -86 0 1 -12620
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_4  sky130_fd_sc_hd__clkinv_4_9
timestamp 1633901636
transform 1 0 -730 0 1 -12620
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_5
timestamp 1633901636
transform 1 0 -2294 0 1 -12620
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_16  sky130_fd_sc_hd__clkbuf_16_5
timestamp 1633901636
transform 1 0 -1926 0 -1 -12620
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_8  sky130_fd_sc_hd__clkbuf_8_4
timestamp 1633901636
transform 1 0 558 0 1 -12620
box -38 -48 1050 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_23
timestamp 1633901636
transform 1 0 -2202 0 1 -12620
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_22
timestamp 1633901636
transform 1 0 -1466 0 1 -12620
box -38 -48 774 592
use n-leg  n-leg_4
timestamp 1643392248
transform 1 0 -284 0 1 -12620
box 1854 -48 6546 1136
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_17
timestamp 1633901636
transform 1 0 -86 0 1 -11532
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_16
timestamp 1633901636
transform 1 0 -86 0 1 -10444
box -38 -48 130 592
use p-leg  p-leg_4
timestamp 1643671812
transform 1 0 2 0 1 -11542
box -34 -38 6666 2234
use sky130_fd_sc_hd__clkinv_16  sky130_fd_sc_hd__clkinv_16_12
timestamp 1633901636
transform 1 0 -2294 0 1 -11532
box -38 -48 2246 592
use sky130_fd_sc_hd__clkinv_16  sky130_fd_sc_hd__clkinv_16_13
timestamp 1633901636
transform 1 0 -2294 0 -1 -10444
box -38 -48 2246 592
use sky130_fd_sc_hd__clkinv_16  sky130_fd_sc_hd__clkinv_16_14
timestamp 1633901636
transform 1 0 -2294 0 1 -10444
box -38 -48 2246 592
use sky130_fd_sc_hd__clkinv_4  sky130_fd_sc_hd__clkinv_4_6
timestamp 1633901636
transform 1 0 -86 0 1 -9356
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_4  sky130_fd_sc_hd__clkinv_4_7
timestamp 1633901636
transform 1 0 -730 0 1 -9356
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_4
timestamp 1633901636
transform 1 0 -2294 0 1 -9356
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_8  sky130_fd_sc_hd__clkbuf_8_3
timestamp 1633901636
transform 1 0 558 0 1 -9356
box -38 -48 1050 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_21
timestamp 1633901636
transform 1 0 -2202 0 1 -9356
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_20
timestamp 1633901636
transform 1 0 -1466 0 1 -9356
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_16  sky130_fd_sc_hd__clkbuf_16_4
timestamp 1633901636
transform 1 0 -1926 0 -1 -9356
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_15
timestamp 1633901636
transform 1 0 -86 0 1 -8268
box -38 -48 130 592
use sky130_fd_sc_hd__clkinv_16  sky130_fd_sc_hd__clkinv_16_9
timestamp 1633901636
transform 1 0 -2294 0 1 -8268
box -38 -48 2246 592
use n-leg  n-leg_3
timestamp 1643392248
transform 1 0 -284 0 1 -9356
box 1854 -48 6546 1136
use p-leg  p-leg_3
timestamp 1643671812
transform 1 0 2 0 1 -8278
box -34 -38 6666 2234
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_14
timestamp 1633901636
transform 1 0 -86 0 1 -7180
box -38 -48 130 592
use sky130_fd_sc_hd__clkinv_16  sky130_fd_sc_hd__clkinv_16_11
timestamp 1633901636
transform 1 0 -2294 0 1 -7180
box -38 -48 2246 592
use sky130_fd_sc_hd__clkinv_16  sky130_fd_sc_hd__clkinv_16_10
timestamp 1633901636
transform 1 0 -2294 0 -1 -7180
box -38 -48 2246 592
use sky130_fd_sc_hd__clkinv_4  sky130_fd_sc_hd__clkinv_4_4
timestamp 1633901636
transform 1 0 -86 0 1 -6092
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_4  sky130_fd_sc_hd__clkinv_4_5
timestamp 1633901636
transform 1 0 -730 0 1 -6092
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_3
timestamp 1633901636
transform 1 0 -2294 0 1 -6092
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_16  sky130_fd_sc_hd__clkbuf_16_3
timestamp 1633901636
transform 1 0 -1926 0 -1 -6092
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_8  sky130_fd_sc_hd__clkbuf_8_2
timestamp 1633901636
transform 1 0 558 0 1 -6092
box -38 -48 1050 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_19
timestamp 1633901636
transform 1 0 -2202 0 1 -6092
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_18
timestamp 1633901636
transform 1 0 -1466 0 1 -6092
box -38 -48 774 592
use n-leg  n-leg_2
timestamp 1643392248
transform 1 0 -284 0 1 -6092
box 1854 -48 6546 1136
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_13
timestamp 1633901636
transform 1 0 -86 0 1 -5004
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_12
timestamp 1633901636
transform 1 0 -86 0 1 -3916
box -38 -48 130 592
use p-leg  p-leg_2
timestamp 1643671812
transform 1 0 2 0 1 -5014
box -34 -38 6666 2234
use sky130_fd_sc_hd__clkinv_16  sky130_fd_sc_hd__clkinv_16_6
timestamp 1633901636
transform 1 0 -2294 0 1 -5004
box -38 -48 2246 592
use sky130_fd_sc_hd__clkinv_16  sky130_fd_sc_hd__clkinv_16_8
timestamp 1633901636
transform 1 0 -2294 0 1 -3916
box -38 -48 2246 592
use sky130_fd_sc_hd__clkinv_16  sky130_fd_sc_hd__clkinv_16_7
timestamp 1633901636
transform 1 0 -2294 0 -1 -3916
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_16  sky130_fd_sc_hd__clkbuf_16_2
timestamp 1633901636
transform 1 0 -1926 0 -1 -2828
box -38 -48 1878 592
use sky130_fd_sc_hd__clkinv_4  sky130_fd_sc_hd__clkinv_4_2
timestamp 1633901636
transform 1 0 -86 0 1 -2828
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_4  sky130_fd_sc_hd__clkinv_4_3
timestamp 1633901636
transform 1 0 -730 0 1 -2828
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_2
timestamp 1633901636
transform 1 0 -2294 0 1 -2828
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_8  sky130_fd_sc_hd__clkbuf_8_1
timestamp 1633901636
transform 1 0 558 0 1 -2828
box -38 -48 1050 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_17
timestamp 1633901636
transform 1 0 -2202 0 1 -2828
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_16
timestamp 1633901636
transform 1 0 -1466 0 1 -2828
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_10
timestamp 1633901636
transform 1 0 -86 0 1 -1740
box -38 -48 130 592
use sky130_fd_sc_hd__clkinv_16  sky130_fd_sc_hd__clkinv_16_3
timestamp 1633901636
transform 1 0 -2294 0 1 -1740
box -38 -48 2246 592
use sky130_fd_sc_hd__clkinv_16  sky130_fd_sc_hd__clkinv_16_4
timestamp 1633901636
transform 1 0 -2294 0 -1 -652
box -38 -48 2246 592
use p-leg  p-leg_1
timestamp 1643671812
transform 1 0 2 0 1 -1750
box -34 -38 6666 2234
use n-leg  n-leg_1
timestamp 1643392248
transform 1 0 -284 0 1 -2828
box 1854 -48 6546 1136
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_11
timestamp 1633901636
transform 1 0 -86 0 1 -652
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_16  sky130_fd_sc_hd__clkbuf_16_1
timestamp 1633901636
transform 1 0 -1926 0 -1 436
box -38 -48 1878 592
use sky130_fd_sc_hd__clkinv_16  sky130_fd_sc_hd__clkinv_16_5
timestamp 1633901636
transform 1 0 -2294 0 1 -652
box -38 -48 2246 592
use sky130_fd_sc_hd__clkinv_4  sky130_fd_sc_hd__clkinv_4_1
timestamp 1633901636
transform 1 0 -730 0 1 436
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_4  sky130_fd_sc_hd__clkinv_4_0
timestamp 1633901636
transform 1 0 -86 0 1 436
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_1
timestamp 1633901636
transform 1 0 -2294 0 1 436
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_8  sky130_fd_sc_hd__clkbuf_8_0
timestamp 1633901636
transform 1 0 558 0 1 436
box -38 -48 1050 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_15
timestamp 1633901636
transform 1 0 -2202 0 1 436
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_14
timestamp 1633901636
transform 1 0 -1466 0 1 436
box -38 -48 774 592
use n-leg  n-leg_0
timestamp 1643392248
transform 1 0 -284 0 1 436
box 1854 -48 6546 1136
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_9
timestamp 1633901636
transform 1 0 -86 0 1 1524
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_8
timestamp 1633901636
transform 1 0 -86 0 1 2612
box -38 -48 130 592
use sky130_fd_sc_hd__clkinv_16  sky130_fd_sc_hd__clkinv_16_0
timestamp 1633901636
transform 1 0 -2294 0 1 1524
box -38 -48 2246 592
use p-leg  p-leg_0
timestamp 1643671812
transform 1 0 2 0 1 1514
box -34 -38 6666 2234
use sky130_fd_sc_hd__clkinv_16  sky130_fd_sc_hd__clkinv_16_1
timestamp 1633901636
transform 1 0 -2294 0 -1 2612
box -38 -48 2246 592
use sky130_fd_sc_hd__clkinv_16  sky130_fd_sc_hd__clkinv_16_2
timestamp 1633901636
transform 1 0 -2294 0 1 2612
box -38 -48 2246 592
use sky130_fd_sc_hd__clkbuf_16  sky130_fd_sc_hd__clkbuf_16_0
timestamp 1633901636
transform 1 0 -1926 0 -1 3700
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_1  sky130_fd_sc_hd__fill_1_0
timestamp 1633901636
transform 1 0 -2294 0 1 3700
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_12
timestamp 1633901636
transform 1 0 -1466 0 1 3700
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_13
timestamp 1633901636
transform 1 0 -2202 0 1 3700
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_11
timestamp 1633901636
transform 1 0 -730 0 1 3700
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_1
timestamp 1633901636
transform 1 0 742 0 1 3700
box -38 -48 774 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1633901636
transform 1 0 742 0 1 3700
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_1
timestamp 1633901636
transform 1 0 466 0 1 3700
box -38 -48 314 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_0
timestamp 1633901636
transform 1 0 6 0 1 3700
box -38 -48 774 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_0
timestamp 1633901636
transform 1 0 190 0 1 3700
box -38 -48 314 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_2
timestamp 1633901636
transform 1 0 1478 0 1 3700
box -38 -48 774 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_3
timestamp 1633901636
transform 1 0 1018 0 1 3700
box -38 -48 314 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_4
timestamp 1633901636
transform 1 0 2950 0 1 3700
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_3
timestamp 1633901636
transform 1 0 2214 0 1 3700
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_5
timestamp 1633901636
transform 1 0 3686 0 1 3700
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_7
timestamp 1633901636
transform 1 0 5158 0 1 3700
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_6
timestamp 1633901636
transform 1 0 4422 0 1 3700
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_8
timestamp 1633901636
transform 1 0 5894 0 1 3700
box -38 -48 774 592
<< labels >>
flabel metal2 3696 -18799 3785 3396 1 FreeSerif 6400 0 0 0 DQ
port 0 n
flabel metal2 s 250 3980 308 4292 1 FreeSerif 480 315 0 0 pu_cal_ctrl[0]
port 13 n
flabel metal2 s 526 3980 584 4292 1 FreeSerif 480 315 0 0 pu_cal_ctrl[1]
port 14 n
flabel metal2 s 801 3980 859 4292 1 FreeSerif 480 315 0 0 pu_cal_ctrl[2]
port 15 n
flabel metal2 s 1076 3980 1134 4292 1 FreeSerif 480 315 0 0 pu_cal_ctrl[3]
port 16 n
flabel metal2 s 1633 3980 1691 4292 1 FreeSerif 480 315 0 0 pd_cal_ctrl[0]
port 2 n
flabel metal2 s 1753 3980 1811 4292 1 FreeSerif 480 315 0 0 pd_cal_ctrl[1]
port 3 n
flabel metal2 s 1873 3980 1931 4292 1 FreeSerif 480 315 0 0 pd_cal_ctrl[2]
port 4 n
flabel metal2 s 1993 3980 2051 4292 1 FreeSerif 480 315 0 0 pd_cal_ctrl[3]
port 5 n
flabel metal1 s -2294 4227 -2265 4261 7 FreeSerif 800 0 0 0 VDD
port 24 n
flabel metal1 s -2294 3683 -2265 3717 7 FreeSerif 800 0 0 0 GND
port 1 n
flabel locali s -1909 3485 -1846 3547 7 FreeSerif 480 0 0 0 pu_ctrl[0]
port 17 w
flabel locali s -641 649 -615 694 7 FreeSerif 480 0 0 0 pd_ctrl[0]
port 6 w
flabel locali s -1909 221 -1846 283 7 FreeSerif 480 0 0 0 pu_ctrl[1]
port 18 w
flabel locali s -1909 -3043 -1846 -2981 7 FreeSerif 480 0 0 0 pu_ctrl[2]
port 19 w
flabel locali s -1909 -6307 -1846 -6245 7 FreeSerif 480 0 0 0 pu_ctrl[3]
port 20 w
flabel locali s -1909 -9571 -1846 -9509 7 FreeSerif 480 0 0 0 pu_ctrl[4]
port 21 w
flabel locali s -1909 -12835 -1846 -12773 7 FreeSerif 480 0 0 0 pu_ctrl[5]
port 22 w
flabel locali s -1909 -16099 -1846 -16037 7 FreeSerif 480 0 0 0 pu_ctrl[6]
port 23 w
flabel locali s -641 -2615 -615 -2570 7 FreeSerif 480 0 0 0 pd_ctrl[1]
port 7 w
flabel locali s -641 -5879 -615 -5834 7 FreeSerif 480 0 0 0 pd_ctrl[2]
port 8 w
flabel locali s -641 -9143 -615 -9098 7 FreeSerif 480 0 0 0 pd_ctrl[3]
port 9 w
flabel locali s -641 -12407 -615 -12362 7 FreeSerif 480 0 0 0 pd_ctrl[4]
port 10 w
flabel locali s -641 -15671 -615 -15626 7 FreeSerif 480 0 0 0 pd_ctrl[5]
port 11 w
flabel locali s -641 -18935 -615 -18890 7 FreeSerif 480 0 0 0 pd_ctrl[6]
port 12 w
<< end >>
