**.subckt sstl_res_tb
vtest DQ VDDQ 0
.save  i(vtest)
X1 DQ pd_ctrl[6] pd_ctrl[5] pd_ctrl[4] pd_ctrl[3] pd_ctrl[2] pd_ctrl[1] pd_ctrl[0] pu_ctrl[6]
+ pu_ctrl[5] pu_ctrl[4] pu_ctrl[3] pu_ctrl[2] pu_ctrl[1] pu_ctrl[0] pd_cal[27] pd_cal[26] pd_cal[25] pd_cal[24]
+ pd_cal[23] pd_cal[22] pd_cal[21] pd_cal[20] pd_cal[19] pd_cal[18] pd_cal[17] pd_cal[16] pd_cal[15] pd_cal[14]
+ pd_cal[13] pd_cal[12] pd_cal[11] pd_cal[10] pd_cal[9] pd_cal[8] pd_cal[7] pd_cal[6] pd_cal[5] pd_cal[4]
+ pd_cal[3] pd_cal[2] pd_cal[1] pd_cal[0] pu_cal[27] pu_cal[26] pu_cal[25] pu_cal[24] pu_cal[23] pu_cal[22]
+ pu_cal[21] pu_cal[20] pu_cal[19] pu_cal[18] pu_cal[17] pu_cal[16] pu_cal[15] pu_cal[14] pu_cal[13] pu_cal[12]
+ pu_cal[11] pu_cal[10] pu_cal[9] pu_cal[8] pu_cal[7] pu_cal[6] pu_cal[5] pu_cal[4] pu_cal[3] pu_cal[2]
+ pu_cal[1] pu_cal[0] SSTL
**** begin user architecture code
 ** Local library links to pdk
.lib ./libs/SED_process_SED_lib.spice SED_process_SED
.include /gro/cad/pdk/sky130A/libs.ref/sky130_fd_sc_hd/spice/sky130_fd_sc_hd.spice

**** end user architecture code
**.ends

* expanding   symbol:  SSTL.sym # of pins=5
* sym_path: /mnt/users/ssd2/homes/hinesd3/proj/sstl-design/SSTL.sym
* sch_path: /mnt/users/ssd2/homes/hinesd3/proj/sstl-design/SSTL.sch
.subckt SSTL  DQ  pd_ctrl[6] pd_ctrl[5] pd_ctrl[4] pd_ctrl[3] pd_ctrl[2] pd_ctrl[1] pd_ctrl[0]
+  pu_ctrl[6] pu_ctrl[5] pu_ctrl[4] pu_ctrl[3] pu_ctrl[2] pu_ctrl[1] pu_ctrl[0]  pd_cal_ctrl[27] pd_cal_ctrl[26]
+ pd_cal_ctrl[25] pd_cal_ctrl[24] pd_cal_ctrl[23] pd_cal_ctrl[22] pd_cal_ctrl[21] pd_cal_ctrl[20] pd_cal_ctrl[19]
+ pd_cal_ctrl[18] pd_cal_ctrl[17] pd_cal_ctrl[16] pd_cal_ctrl[15] pd_cal_ctrl[14] pd_cal_ctrl[13] pd_cal_ctrl[12]
+ pd_cal_ctrl[11] pd_cal_ctrl[10] pd_cal_ctrl[9] pd_cal_ctrl[8] pd_cal_ctrl[7] pd_cal_ctrl[6] pd_cal_ctrl[5]
+ pd_cal_ctrl[4] pd_cal_ctrl[3] pd_cal_ctrl[2] pd_cal_ctrl[1] pd_cal_ctrl[0]  pu_cal_ctrl[27] pu_cal_ctrl[26]
+ pu_cal_ctrl[25] pu_cal_ctrl[24] pu_cal_ctrl[23] pu_cal_ctrl[22] pu_cal_ctrl[21] pu_cal_ctrl[20] pu_cal_ctrl[19]
+ pu_cal_ctrl[18] pu_cal_ctrl[17] pu_cal_ctrl[16] pu_cal_ctrl[15] pu_cal_ctrl[14] pu_cal_ctrl[13] pu_cal_ctrl[12]
+ pu_cal_ctrl[11] pu_cal_ctrl[10] pu_cal_ctrl[9] pu_cal_ctrl[8] pu_cal_ctrl[7] pu_cal_ctrl[6] pu_cal_ctrl[5]
+ pu_cal_ctrl[4] pu_cal_ctrl[3] pu_cal_ctrl[2] pu_cal_ctrl[1] pu_cal_ctrl[0]
*.iopin DQ
*.ipin
*+ pu_cal_ctrl[27],pu_cal_ctrl[26],pu_cal_ctrl[25],pu_cal_ctrl[24],pu_cal_ctrl[23],pu_cal_ctrl[22],pu_cal_ctrl[21],pu_cal_ctrl[20],pu_cal_ctrl[19],pu_cal_ctrl[18],pu_cal_ctrl[17],pu_cal_ctrl[16],pu_cal_ctrl[15],pu_cal_ctrl[14],pu_cal_ctrl[13],pu_cal_ctrl[12],pu_cal_ctrl[11],pu_cal_ctrl[10],pu_cal_ctrl[9],pu_cal_ctrl[8],pu_cal_ctrl[7],pu_cal_ctrl[6],pu_cal_ctrl[5],pu_cal_ctrl[4],pu_cal_ctrl[3],pu_cal_ctrl[2],pu_cal_ctrl[1],pu_cal_ctrl[0]
*.ipin
*+ pd_cal_ctrl[27],pd_cal_ctrl[26],pd_cal_ctrl[25],pd_cal_ctrl[24],pd_cal_ctrl[23],pd_cal_ctrl[22],pd_cal_ctrl[21],pd_cal_ctrl[20],pd_cal_ctrl[19],pd_cal_ctrl[18],pd_cal_ctrl[17],pd_cal_ctrl[16],pd_cal_ctrl[15],pd_cal_ctrl[14],pd_cal_ctrl[13],pd_cal_ctrl[12],pd_cal_ctrl[11],pd_cal_ctrl[10],pd_cal_ctrl[9],pd_cal_ctrl[8],pd_cal_ctrl[7],pd_cal_ctrl[6],pd_cal_ctrl[5],pd_cal_ctrl[4],pd_cal_ctrl[3],pd_cal_ctrl[2],pd_cal_ctrl[1],pd_cal_ctrl[0]
*.ipin pu_ctrl[6],pu_ctrl[5],pu_ctrl[4],pu_ctrl[3],pu_ctrl[2],pu_ctrl[1],pu_ctrl[0]
*.ipin pd_ctrl[6],pd_ctrl[5],pd_ctrl[4],pd_ctrl[3],pd_ctrl[2],pd_ctrl[1],pd_ctrl[0]
X1 DQ n_pu_ctrl[6] n_pu_cal_ctrl[27] n_pu_cal_ctrl[26] n_pu_cal_ctrl[25] n_pu_cal_ctrl[24] p-leg
X2 DQ pd_ctrl[6] pd_cal_ctrl[27] pd_cal_ctrl[26] pd_cal_ctrl[25] pd_cal_ctrl[24] n-leg
X3 DQ n_pu_ctrl[5] n_pu_cal_ctrl[23] n_pu_cal_ctrl[22] n_pu_cal_ctrl[21] n_pu_cal_ctrl[20] p-leg
X4 DQ pd_ctrl[5] pd_cal_ctrl[23] pd_cal_ctrl[22] pd_cal_ctrl[21] pd_cal_ctrl[20] n-leg
X5 DQ n_pu_ctrl[4] n_pu_cal_ctrl[19] n_pu_cal_ctrl[18] n_pu_cal_ctrl[17] n_pu_cal_ctrl[16] p-leg
X6 DQ pd_ctrl[4] pd_cal_ctrl[19] pd_cal_ctrl[18] pd_cal_ctrl[17] pd_cal_ctrl[16] n-leg
X7 DQ n_pu_ctrl[3] n_pu_cal_ctrl[15] n_pu_cal_ctrl[14] n_pu_cal_ctrl[13] n_pu_cal_ctrl[12] p-leg
X8 DQ pd_ctrl[3] pd_cal_ctrl[15] pd_cal_ctrl[14] pd_cal_ctrl[13] pd_cal_ctrl[12] n-leg
X9 DQ n_pu_ctrl[2] n_pu_cal_ctrl[11] n_pu_cal_ctrl[10] n_pu_cal_ctrl[9] n_pu_cal_ctrl[8] p-leg
X10 DQ pd_ctrl[2] pd_cal_ctrl[11] pd_cal_ctrl[10] pd_cal_ctrl[9] pd_cal_ctrl[8] n-leg
X11 DQ n_pu_ctrl[1] n_pu_cal_ctrl[7] n_pu_cal_ctrl[6] n_pu_cal_ctrl[5] n_pu_cal_ctrl[4] p-leg
X12 DQ pd_ctrl[1] pd_cal_ctrl[7] pd_cal_ctrl[6] pd_cal_ctrl[5] pd_cal_ctrl[4] n-leg
X13 DQ n_pu_ctrl[0] n_pu_cal_ctrl[3] n_pu_cal_ctrl[2] n_pu_cal_ctrl[1] n_pu_cal_ctrl[0] p-leg
X14 DQ pd_ctrl[0] pd_cal_ctrl[3] pd_cal_ctrl[2] pd_cal_ctrl[1] pd_cal_ctrl[0] n-leg
xpd_buff_4[6] pd_ctrl[6] VGND VNB VPB VPWR pdc4[6] sky130_fd_sc_hd__inv_4
xpd_buff_4[5] pd_ctrl[5] VGND VNB VPB VPWR pdc4[5] sky130_fd_sc_hd__inv_4
xpd_buff_4[4] pd_ctrl[4] VGND VNB VPB VPWR pdc4[4] sky130_fd_sc_hd__inv_4
xpd_buff_4[3] pd_ctrl[3] VGND VNB VPB VPWR pdc4[3] sky130_fd_sc_hd__inv_4
xpd_buff_4[2] pd_ctrl[2] VGND VNB VPB VPWR pdc4[2] sky130_fd_sc_hd__inv_4
xpd_buff_4[1] pd_ctrl[1] VGND VNB VPB VPWR pdc4[1] sky130_fd_sc_hd__inv_4
xpd_buff_4[0] pd_ctrl[0] VGND VNB VPB VPWR pdc4[0] sky130_fd_sc_hd__inv_4
xpd_buff_6[6] pdc4[6] VGND VNB VPB VPWR pd_ctrl[6] sky130_fd_sc_hd__inv_6
xpd_buff_6[5] pdc4[5] VGND VNB VPB VPWR pd_ctrl[5] sky130_fd_sc_hd__inv_6
xpd_buff_6[4] pdc4[4] VGND VNB VPB VPWR pd_ctrl[4] sky130_fd_sc_hd__inv_6
xpd_buff_6[3] pdc4[3] VGND VNB VPB VPWR pd_ctrl[3] sky130_fd_sc_hd__inv_6
xpd_buff_6[2] pdc4[2] VGND VNB VPB VPWR pd_ctrl[2] sky130_fd_sc_hd__inv_6
xpd_buff_6[1] pdc4[1] VGND VNB VPB VPWR pd_ctrl[1] sky130_fd_sc_hd__inv_6
xpd_buff_6[0] pdc4[0] VGND VNB VPB VPWR pd_ctrl[0] sky130_fd_sc_hd__inv_6
xpu_buff_4[6] puc1[6] VGND VNB VPB VPWR puc4[6] sky130_fd_sc_hd__inv_4
xpu_buff_4[5] puc1[5] VGND VNB VPB VPWR puc4[5] sky130_fd_sc_hd__inv_4
xpu_buff_4[4] puc1[4] VGND VNB VPB VPWR puc4[4] sky130_fd_sc_hd__inv_4
xpu_buff_4[3] puc1[3] VGND VNB VPB VPWR puc4[3] sky130_fd_sc_hd__inv_4
xpu_buff_4[2] puc1[2] VGND VNB VPB VPWR puc4[2] sky130_fd_sc_hd__inv_4
xpu_buff_4[1] puc1[1] VGND VNB VPB VPWR puc4[1] sky130_fd_sc_hd__inv_4
xpu_buff_4[0] puc1[0] VGND VNB VPB VPWR puc4[0] sky130_fd_sc_hd__inv_4
xpu_buff_6[6] puc4[6] VGND VNB VPB VPWR n_pu_ctrl[6] sky130_fd_sc_hd__inv_6
xpu_buff_6[5] puc4[5] VGND VNB VPB VPWR n_pu_ctrl[5] sky130_fd_sc_hd__inv_6
xpu_buff_6[4] puc4[4] VGND VNB VPB VPWR n_pu_ctrl[4] sky130_fd_sc_hd__inv_6
xpu_buff_6[3] puc4[3] VGND VNB VPB VPWR n_pu_ctrl[3] sky130_fd_sc_hd__inv_6
xpu_buff_6[2] puc4[2] VGND VNB VPB VPWR n_pu_ctrl[2] sky130_fd_sc_hd__inv_6
xpu_buff_6[1] puc4[1] VGND VNB VPB VPWR n_pu_ctrl[1] sky130_fd_sc_hd__inv_6
xpu_buff_6[0] puc4[0] VGND VNB VPB VPWR n_pu_ctrl[0] sky130_fd_sc_hd__inv_6
xpu_buff_1[6] pu_ctrl[6] VGND VNB VPB VPWR puc1[6] sky130_fd_sc_hd__inv_1
xpu_buff_1[5] pu_ctrl[5] VGND VNB VPB VPWR puc1[5] sky130_fd_sc_hd__inv_1
xpu_buff_1[4] pu_ctrl[4] VGND VNB VPB VPWR puc1[4] sky130_fd_sc_hd__inv_1
xpu_buff_1[3] pu_ctrl[3] VGND VNB VPB VPWR puc1[3] sky130_fd_sc_hd__inv_1
xpu_buff_1[2] pu_ctrl[2] VGND VNB VPB VPWR puc1[2] sky130_fd_sc_hd__inv_1
xpu_buff_1[1] pu_ctrl[1] VGND VNB VPB VPWR puc1[1] sky130_fd_sc_hd__inv_1
xpu_buff_1[0] pu_ctrl[0] VGND VNB VPB VPWR puc1[0] sky130_fd_sc_hd__inv_1
xpu_cal_inv[27] pu_cal_ctrl[27] VGND VNB VPB VPWR n_pu_cal_ctrl[27] sky130_fd_sc_hd__inv_1
xpu_cal_inv[26] pu_cal_ctrl[26] VGND VNB VPB VPWR n_pu_cal_ctrl[26] sky130_fd_sc_hd__inv_1
xpu_cal_inv[25] pu_cal_ctrl[25] VGND VNB VPB VPWR n_pu_cal_ctrl[25] sky130_fd_sc_hd__inv_1
xpu_cal_inv[24] pu_cal_ctrl[24] VGND VNB VPB VPWR n_pu_cal_ctrl[24] sky130_fd_sc_hd__inv_1
xpu_cal_inv[23] pu_cal_ctrl[23] VGND VNB VPB VPWR n_pu_cal_ctrl[23] sky130_fd_sc_hd__inv_1
xpu_cal_inv[22] pu_cal_ctrl[22] VGND VNB VPB VPWR n_pu_cal_ctrl[22] sky130_fd_sc_hd__inv_1
xpu_cal_inv[21] pu_cal_ctrl[21] VGND VNB VPB VPWR n_pu_cal_ctrl[21] sky130_fd_sc_hd__inv_1
xpu_cal_inv[20] pu_cal_ctrl[20] VGND VNB VPB VPWR n_pu_cal_ctrl[20] sky130_fd_sc_hd__inv_1
xpu_cal_inv[19] pu_cal_ctrl[19] VGND VNB VPB VPWR n_pu_cal_ctrl[19] sky130_fd_sc_hd__inv_1
xpu_cal_inv[18] pu_cal_ctrl[18] VGND VNB VPB VPWR n_pu_cal_ctrl[18] sky130_fd_sc_hd__inv_1
xpu_cal_inv[17] pu_cal_ctrl[17] VGND VNB VPB VPWR n_pu_cal_ctrl[17] sky130_fd_sc_hd__inv_1
xpu_cal_inv[16] pu_cal_ctrl[16] VGND VNB VPB VPWR n_pu_cal_ctrl[16] sky130_fd_sc_hd__inv_1
xpu_cal_inv[15] pu_cal_ctrl[15] VGND VNB VPB VPWR n_pu_cal_ctrl[15] sky130_fd_sc_hd__inv_1
xpu_cal_inv[14] pu_cal_ctrl[14] VGND VNB VPB VPWR n_pu_cal_ctrl[14] sky130_fd_sc_hd__inv_1
xpu_cal_inv[13] pu_cal_ctrl[13] VGND VNB VPB VPWR n_pu_cal_ctrl[13] sky130_fd_sc_hd__inv_1
xpu_cal_inv[12] pu_cal_ctrl[12] VGND VNB VPB VPWR n_pu_cal_ctrl[12] sky130_fd_sc_hd__inv_1
xpu_cal_inv[11] pu_cal_ctrl[11] VGND VNB VPB VPWR n_pu_cal_ctrl[11] sky130_fd_sc_hd__inv_1
xpu_cal_inv[10] pu_cal_ctrl[10] VGND VNB VPB VPWR n_pu_cal_ctrl[10] sky130_fd_sc_hd__inv_1
xpu_cal_inv[9] pu_cal_ctrl[9] VGND VNB VPB VPWR n_pu_cal_ctrl[9] sky130_fd_sc_hd__inv_1
xpu_cal_inv[8] pu_cal_ctrl[8] VGND VNB VPB VPWR n_pu_cal_ctrl[8] sky130_fd_sc_hd__inv_1
xpu_cal_inv[7] pu_cal_ctrl[7] VGND VNB VPB VPWR n_pu_cal_ctrl[7] sky130_fd_sc_hd__inv_1
xpu_cal_inv[6] pu_cal_ctrl[6] VGND VNB VPB VPWR n_pu_cal_ctrl[6] sky130_fd_sc_hd__inv_1
xpu_cal_inv[5] pu_cal_ctrl[5] VGND VNB VPB VPWR n_pu_cal_ctrl[5] sky130_fd_sc_hd__inv_1
xpu_cal_inv[4] pu_cal_ctrl[4] VGND VNB VPB VPWR n_pu_cal_ctrl[4] sky130_fd_sc_hd__inv_1
xpu_cal_inv[3] pu_cal_ctrl[3] VGND VNB VPB VPWR n_pu_cal_ctrl[3] sky130_fd_sc_hd__inv_1
xpu_cal_inv[2] pu_cal_ctrl[2] VGND VNB VPB VPWR n_pu_cal_ctrl[2] sky130_fd_sc_hd__inv_1
xpu_cal_inv[1] pu_cal_ctrl[1] VGND VNB VPB VPWR n_pu_cal_ctrl[1] sky130_fd_sc_hd__inv_1
xpu_cal_inv[0] pu_cal_ctrl[0] VGND VNB VPB VPWR n_pu_cal_ctrl[0] sky130_fd_sc_hd__inv_1
V1 VDD VPWR 0
V2 VGND GND 0
V3 VDD VPB 0
V4 VNB GND 0
.ends


* expanding   symbol:  p-leg.sym # of pins=3
* sym_path: /mnt/users/ssd2/homes/hinesd3/proj/sstl-design/p-leg.sym
* sch_path: /mnt/users/ssd2/homes/hinesd3/proj/sstl-design/p-leg.sch
.subckt p-leg  DQ  n_pu_ctrl  n_cal_ctrl[3] n_cal_ctrl[2] n_cal_ctrl[1] n_cal_ctrl[0]
*.ipin n_cal_ctrl[3],n_cal_ctrl[2],n_cal_ctrl[1],n_cal_ctrl[0]
*.ipin n_pu_ctrl
*.iopin DQ
R1 DQ net1 sky130_fd_pr__res_generic_po W=0.33 L=1.8 m=1
XMpullup net1 n_pu_ctrl VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=128 m=128
XMctrltot VDD n_cal_ctrl[0] VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=120 m=120
XMctrl0 DQ n_cal_ctrl[0] net1 VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=48 m=48
XMctrl1 DQ n_cal_ctrl[1] net1 VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=16 m=16
XMctrl2 DQ n_cal_ctrl[2] net1 VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=8 m=8
XMctrl3 DQ n_cal_ctrl[3] net1 VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=4 m=4
.ends


* expanding   symbol:  n-leg.sym # of pins=3
* sym_path: /mnt/users/ssd2/homes/hinesd3/proj/sstl-design/n-leg.sym
* sch_path: /mnt/users/ssd2/homes/hinesd3/proj/sstl-design/n-leg.sch
.subckt n-leg  DQ  pd_ctrl  cal_ctrl[3] cal_ctrl[2] cal_ctrl[1] cal_ctrl[0]
*.iopin DQ
*.ipin pd_ctrl
*.ipin cal_ctrl[3],cal_ctrl[2],cal_ctrl[1],cal_ctrl[0]
R1 vpulldown DQ sky130_fd_pr__res_generic_po W=0.33 L=1.7 m=1
Xn1 vpulldown pd_ctrl GND GND sky130_fd_pr__nfet_01v8 L=0.15 W=0.65 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=48 m=48
Xnctrl0 DQ cal_ctrl[0] vpulldown GND sky130_fd_pr__nfet_01v8 L=0.15 W=0.65 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=6 m=6
Xnctrl1 DQ cal_ctrl[1] vpulldown GND sky130_fd_pr__nfet_01v8 L=0.15 W=0.65 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=3 m=3
Xnctrl2 DQ cal_ctrl[2] vpulldown GND sky130_fd_pr__nfet_01v8 L=0.15 W=0.975 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
Xnctrl3 DQ cal_ctrl[3] vpulldown GND sky130_fd_pr__nfet_01v8 L=0.15 W=0.5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
Xnctrl_tot GND GND GND GND sky130_fd_pr__nfet_01v8 L=0.15 W=0.65 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=11 m=11
.ends

.GLOBAL VDD
.GLOBAL GND
**** begin user architecture code


* power voltage
vvddq VDDQ 0 0
vvdd VDD 0 SED_vdd_SED

** CALIBRATION CONTROL **
* PULLUP
vpu_cal00 pu_cal[0] 0 SED_pucal00_SED
vpu_cal01 pu_cal[1] 0 SED_pucal01_SED
vpu_cal02 pu_cal[2] 0 SED_pucal02_SED
vpu_cal03 pu_cal[3] 0 SED_pucal03_SED
vpu_cal10 pu_cal[4] 0 SED_pucal10_SED
vpu_cal11 pu_cal[5] 0 SED_pucal11_SED
vpu_cal12 pu_cal[6] 0 SED_pucal12_SED
vpu_cal13 pu_cal[7] 0 SED_pucal13_SED
vpu_cal20 pu_cal[8] 0 SED_pucal20_SED
vpu_cal21 pu_cal[9] 0 SED_pucal21_SED
vpu_cal22 pu_cal[10] 0 SED_pucal22_SED
vpu_cal23 pu_cal[11] 0 SED_pucal23_SED
vpu_cal30 pu_cal[12] 0 SED_pucal30_SED
vpu_cal31 pu_cal[13] 0 SED_pucal31_SED
vpu_cal32 pu_cal[14] 0 SED_pucal32_SED
vpu_cal33 pu_cal[15] 0 SED_pucal33_SED
vpu_cal40 pu_cal[16] 0 SED_pucal40_SED
vpu_cal41 pu_cal[17] 0 SED_pucal41_SED
vpu_cal42 pu_cal[18] 0 SED_pucal42_SED
vpu_cal43 pu_cal[19] 0 SED_pucal43_SED
vpu_cal50 pu_cal[20] 0 SED_pucal50_SED
vpu_cal51 pu_cal[21] 0 SED_pucal51_SED
vpu_cal52 pu_cal[22] 0 SED_pucal52_SED
vpu_cal53 pu_cal[23] 0 SED_pucal53_SED
vpu_cal60 pu_cal[24] 0 SED_pucal60_SED
vpu_cal61 pu_cal[25] 0 SED_pucal61_SED
vpu_cal62 pu_cal[26] 0 SED_pucal62_SED
vpu_cal63 pu_cal[27] 0 SED_pucal63_SED
* PULLDOWN
vpd_cal00 pd_cal[0] 0 SED_pdcal00_SED
vpd_cal01 pd_cal[1] 0 SED_pdcal01_SED
vpd_cal02 pd_cal[2] 0 SED_pdcal02_SED
vpd_cal03 pd_cal[3] 0 SED_pdcal03_SED
vpd_cal10 pd_cal[4] 0 SED_pdcal10_SED
vpd_cal11 pd_cal[5] 0 SED_pdcal11_SED
vpd_cal12 pd_cal[6] 0 SED_pdcal12_SED
vpd_cal13 pd_cal[7] 0 SED_pdcal13_SED
vpd_cal20 pd_cal[8] 0 SED_pdcal20_SED
vpd_cal21 pd_cal[9] 0 SED_pdcal21_SED
vpd_cal22 pd_cal[10] 0 SED_pdcal22_SED
vpd_cal23 pd_cal[11] 0 SED_pdcal23_SED
vpd_cal30 pd_cal[12] 0 SED_pdcal30_SED
vpd_cal31 pd_cal[13] 0 SED_pdcal31_SED
vpd_cal32 pd_cal[14] 0 SED_pdcal32_SED
vpd_cal33 pd_cal[15] 0 SED_pdcal33_SED
vpd_cal40 pd_cal[16] 0 SED_pdcal40_SED
vpd_cal41 pd_cal[17] 0 SED_pdcal41_SED
vpd_cal42 pd_cal[18] 0 SED_pdcal42_SED
vpd_cal43 pd_cal[19] 0 SED_pdcal43_SED
vpd_cal50 pd_cal[20] 0 SED_pdcal50_SED
vpd_cal51 pd_cal[21] 0 SED_pdcal51_SED
vpd_cal52 pd_cal[22] 0 SED_pdcal52_SED
vpd_cal53 pd_cal[23] 0 SED_pdcal53_SED
vpd_cal60 pd_cal[24] 0 SED_pdcal60_SED
vpd_cal61 pd_cal[25] 0 SED_pdcal61_SED
vpd_cal62 pd_cal[26] 0 SED_pdcal62_SED
vpd_cal63 pd_cal[27] 0 SED_pdcal63_SED

** LEG ENABLE/DISABLE CONTROL
* PULLUP
vpu_ctrl0 pu_ctrl[0] 0 SED_puctrl0_SED
vpu_ctrl1 pu_ctrl[1] 0 SED_puctrl1_SED
vpu_ctrl2 pu_ctrl[2] 0 SED_puctrl2_SED
vpu_ctrl3 pu_ctrl[3] 0 SED_puctrl3_SED
vpu_ctrl4 pu_ctrl[4] 0 SED_puctrl4_SED
vpu_ctrl5 pu_ctrl[5] 0 SED_puctrl5_SED
vpu_ctrl6 pu_ctrl[6] 0 SED_puctrl6_SED
* PULLDOWN
vpd_ctrl0 pd_ctrl[0] 0 SED_pdctrl0_SED
vpd_ctrl1 pd_ctrl[1] 0 SED_pdctrl1_SED
vpd_ctrl2 pd_ctrl[2] 0 SED_pdctrl2_SED
vpd_ctrl3 pd_ctrl[3] 0 SED_pdctrl3_SED
vpd_ctrl4 pd_ctrl[4] 0 SED_pdctrl4_SED
vpd_ctrl5 pd_ctrl[5] 0 SED_pdctrl5_SED
vpd_ctrl6 pd_ctrl[6] 0 SED_pdctrl6_SED


.control
save all
set temp=SED_temp_SED

* RUN SIMULATION
dc vvddq 0.3 1.2 0.05
* OUTPUT
print v(vddq)/i(vtest)
wrdata out/data/SED_plotName_SED.txt v(vddq)/i(vtest)
set hcopydevtype = svg
hardcopy ./out/plots/SED_plotName_SED.svg vddq/I(vtest) vs vddq title 'Resistance vs pin voltage'

.endc


**** end user architecture code
.end
