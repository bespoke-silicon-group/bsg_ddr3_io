**.subckt test_pu_res
Vgate VDD net1 SED_vg_SED
R1 net3 net2 sky130_fd_pr__res_generic_po W=0.33 L=1.8 m=1
vtest net3 VDDQ 0
.save  i(vtest)
XM2 net4 net4 net4 net4 sky130_fd_pr__pfet_01v8_hvt L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=256 m=256
V1v5 v1v5 GND SED_v1v5_SED
Vpinvoltage v1v5 VDDQ 0
XM1 net5 net5 net5 net5 sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=256 m=256
XM3 net2 net1 v1v5 VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=128 m=128
**** begin user architecture code
 ** Local library links to pdk
.lib ./libs/SED_process_SED_lib.spice SED_process_SED

**** end user architecture code
**.ends
.GLOBAL VDD
.GLOBAL GND
**** begin user architecture code



* power voltage
vvdd VDD 0 1.8

*.param rwidth=4.6

.control
save all
set temp=SED_temp_SED

* RUN SIMULATION
dc Vpinvoltage 0.3 1.2 0.05
* OUTPUT
print (SED_v1v5_SED-vddq)/i(vtest)
wrdata out/data/SED_plotName_SED.txt (SED_v1v5_SED-vddq)/i(vtest)
set hcopydevtype = svg
hardcopy ./out/plots/SED_plotName_SED.svg (SED_v1v5_SED-vddq)/I(vtest) vs vddq title 'Resistance vs pin voltage'

.endc


**** end user architecture code
.end
