**.subckt test_resistance
R1 vpulldown net1 sky130_fd_pr__res_generic_po W=0.33 L=1.73 m=1
vtest VDDQ net1 0
.save  i(vtest)
Xn1 vpulldown net2 GND GND sky130_fd_pr__nfet_01v8 L=0.15 W=0.65 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=64 m=64 
Vgate net2 GND SED_vg_SED
**** begin user architecture code
 ** Local library links to pdk
.lib ./libs/SED_process_SED_lib.spice SED_process_SED

**** end user architecture code
**.ends
.GLOBAL GND
**** begin user architecture code



* power voltage
vvddq VDDQ 0 0
*.param rwidth=4.6

.control
save all
set temp=SED_temp_SED

* RUN SIMULATION
dc vvddq 0.1 1.65 0.05
* OUTPUT
*plot vddq/I(vtest) vs vddq
*MEAS DC r_max MAX par('vddq/I(vtest)')
print v(vddq)/i(vtest)
set hcopydevtype = svg
hardcopy ./out/plots/SED_plotName_SED.svg vddq/I(vtest) vs vddq title 'Resistance vs pin voltage'

.endc


**** end user architecture code
.end
