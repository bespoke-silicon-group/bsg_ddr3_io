* Slow-Fast corner with mismatch (sf_mm)
.lib sf_mm
.param mc_mm_switch=1
.param mc_pr_switch=0
* MOSFET
.include "../../pdk/libs.tech/ngspice/corners/sf.spice"
* Resistor/Capacitor
.include "../../pdk/libs.tech/ngspice/r+c/res_typical__cap_typical.spice"
.include "../../pdk/libs.tech/ngspice/r+c/res_typical__cap_typical__lin.spice"
* Special cells
.include "../../pdk/libs.tech/ngspice/corners/sf/specialized_cells.spice"
.endl sf_mm
