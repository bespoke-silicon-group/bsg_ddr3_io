* High-High corner with mismatch (hh_mm)
.lib hh_mm
.param mc_mm_switch=1
.param mc_pr_switch=0
* MOSFET
.include "sky130_libs/corners/tt.spice"
* Resistor/Capacitor
.include "sky130_libs/r+c/res_high__cap_high.spice"
.include "sky130_libs/r+c/res_high__cap_high__lin.spice"
* Special cells
.include "sky130_libs/corners/tt/specialized_cells.spice"
.endl hh_mm
