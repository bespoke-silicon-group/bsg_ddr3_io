* High-Low corner with mismatch (hl_mm)
.lib hl_mm
.param mc_mm_switch=1
.param mc_pr_switch=0
* MOSFET
.include "../../pdk/libs.tech/ngspice/corners/tt.spice"
* Resistor/Capacitor
.include "../../pdk/libs.tech/ngspice/r+c/res_high__cap_low.spice"
.include "../../pdk/libs.tech/ngspice/r+c/res_high__cap_low__lin.spice"
* Special cells
.include "../../pdk/libs.tech/ngspice/corners/tt/specialized_cells.spice"
.endl hl_mm
