magic
tech sky130A
magscale 1 2
timestamp 1643248389
<< nwell >>
rect -34 1604 6666 1925
rect 6498 271 6666 592
<< pwell >>
rect 30 2162 74 2196
rect 766 2162 810 2196
rect 1501 2162 1545 2196
rect 2237 2162 2281 2196
rect 2973 2162 3017 2196
rect 3709 2162 3753 2196
rect 4445 2162 4489 2196
rect 5181 2162 5225 2196
rect 5917 2162 5961 2196
<< nsubdiff >>
rect 6289 1857 6323 1881
rect 6289 1773 6323 1823
rect 6289 1706 6323 1739
rect 6565 457 6599 490
rect 6565 373 6599 423
rect 6565 315 6599 339
<< nsubdiffcont >>
rect 6289 1823 6323 1857
rect 6289 1739 6323 1773
rect 6565 423 6599 457
rect 6565 339 6599 373
<< poly >>
rect 773 1494 831 1576
rect 1541 1494 1599 1576
rect 2309 1494 2367 1576
rect 4567 1420 4625 1502
<< locali >>
rect 4 2169 33 2203
rect 67 2169 125 2203
rect 159 2169 217 2203
rect 251 2169 309 2203
rect 343 2169 401 2203
rect 435 2169 493 2203
rect 527 2169 585 2203
rect 619 2169 677 2203
rect 711 2169 769 2203
rect 803 2169 861 2203
rect 895 2169 953 2203
rect 987 2169 1045 2203
rect 1079 2169 1137 2203
rect 1171 2169 1229 2203
rect 1263 2169 1321 2203
rect 1355 2169 1413 2203
rect 1447 2169 1504 2203
rect 1538 2169 1596 2203
rect 1630 2169 1688 2203
rect 1722 2169 1780 2203
rect 1814 2169 1872 2203
rect 1906 2169 1964 2203
rect 1998 2169 2056 2203
rect 2090 2169 2148 2203
rect 2182 2169 2240 2203
rect 2274 2169 2332 2203
rect 2366 2169 2424 2203
rect 2458 2169 2516 2203
rect 2550 2169 2608 2203
rect 2642 2169 2700 2203
rect 2734 2169 2792 2203
rect 2826 2169 2884 2203
rect 2918 2169 2976 2203
rect 3010 2169 3068 2203
rect 3102 2169 3160 2203
rect 3194 2169 3252 2203
rect 3286 2169 3344 2203
rect 3378 2169 3436 2203
rect 3470 2169 3528 2203
rect 3562 2169 3620 2203
rect 3654 2169 3712 2203
rect 3746 2169 3804 2203
rect 3838 2169 3896 2203
rect 3930 2169 3988 2203
rect 4022 2169 4080 2203
rect 4114 2169 4172 2203
rect 4206 2169 4264 2203
rect 4298 2169 4356 2203
rect 4390 2169 4448 2203
rect 4482 2169 4540 2203
rect 4574 2169 4632 2203
rect 4666 2169 4724 2203
rect 4758 2169 4816 2203
rect 4850 2169 4908 2203
rect 4942 2169 5000 2203
rect 5034 2169 5092 2203
rect 5126 2169 5184 2203
rect 5218 2169 5276 2203
rect 5310 2169 5368 2203
rect 5402 2169 5460 2203
rect 5494 2169 5552 2203
rect 5586 2169 5644 2203
rect 5678 2169 5736 2203
rect 5770 2169 5828 2203
rect 5862 2169 5920 2203
rect 5954 2169 6012 2203
rect 6046 2169 6104 2203
rect 6138 2169 6196 2203
rect 6230 2169 6288 2203
rect 6322 2169 6380 2203
rect 6414 2169 6472 2203
rect 6506 2169 6564 2203
rect 6598 2169 6628 2203
rect 16 1957 3260 2067
rect 3330 1957 6194 2067
rect 6277 1857 6335 1892
rect 6277 1823 6289 1857
rect 6323 1823 6335 1857
rect 6277 1773 6335 1823
rect 6277 1739 6289 1773
rect 6323 1739 6335 1773
rect 6277 1659 6335 1739
rect 6260 1625 6289 1659
rect 6323 1625 6352 1659
rect 5369 1537 6273 1591
rect 3135 1480 3823 1483
rect 3135 1424 3260 1480
rect 3330 1424 3823 1480
rect 3135 1412 3823 1424
rect 3752 1338 3823 1412
rect 5369 1338 5409 1537
rect 17 1304 3718 1329
rect 17 1264 3845 1304
rect 3594 1255 3845 1264
rect 5443 1255 5483 1454
rect 3594 1248 5483 1255
rect 3718 1164 5483 1248
rect 6536 537 6565 571
rect 6599 537 6628 571
rect 6553 457 6611 537
rect 6553 423 6565 457
rect 6599 423 6611 457
rect 6553 373 6611 423
rect 6553 339 6565 373
rect 6599 339 6611 373
rect 6553 304 6611 339
<< viali >>
rect 33 2169 67 2203
rect 125 2169 159 2203
rect 217 2169 251 2203
rect 309 2169 343 2203
rect 401 2169 435 2203
rect 493 2169 527 2203
rect 585 2169 619 2203
rect 677 2169 711 2203
rect 769 2169 803 2203
rect 861 2169 895 2203
rect 953 2169 987 2203
rect 1045 2169 1079 2203
rect 1137 2169 1171 2203
rect 1229 2169 1263 2203
rect 1321 2169 1355 2203
rect 1413 2169 1447 2203
rect 1504 2169 1538 2203
rect 1596 2169 1630 2203
rect 1688 2169 1722 2203
rect 1780 2169 1814 2203
rect 1872 2169 1906 2203
rect 1964 2169 1998 2203
rect 2056 2169 2090 2203
rect 2148 2169 2182 2203
rect 2240 2169 2274 2203
rect 2332 2169 2366 2203
rect 2424 2169 2458 2203
rect 2516 2169 2550 2203
rect 2608 2169 2642 2203
rect 2700 2169 2734 2203
rect 2792 2169 2826 2203
rect 2884 2169 2918 2203
rect 2976 2169 3010 2203
rect 3068 2169 3102 2203
rect 3160 2169 3194 2203
rect 3252 2169 3286 2203
rect 3344 2169 3378 2203
rect 3436 2169 3470 2203
rect 3528 2169 3562 2203
rect 3620 2169 3654 2203
rect 3712 2169 3746 2203
rect 3804 2169 3838 2203
rect 3896 2169 3930 2203
rect 3988 2169 4022 2203
rect 4080 2169 4114 2203
rect 4172 2169 4206 2203
rect 4264 2169 4298 2203
rect 4356 2169 4390 2203
rect 4448 2169 4482 2203
rect 4540 2169 4574 2203
rect 4632 2169 4666 2203
rect 4724 2169 4758 2203
rect 4816 2169 4850 2203
rect 4908 2169 4942 2203
rect 5000 2169 5034 2203
rect 5092 2169 5126 2203
rect 5184 2169 5218 2203
rect 5276 2169 5310 2203
rect 5368 2169 5402 2203
rect 5460 2169 5494 2203
rect 5552 2169 5586 2203
rect 5644 2169 5678 2203
rect 5736 2169 5770 2203
rect 5828 2169 5862 2203
rect 5920 2169 5954 2203
rect 6012 2169 6046 2203
rect 6104 2169 6138 2203
rect 6196 2169 6230 2203
rect 6288 2169 6322 2203
rect 6380 2169 6414 2203
rect 6472 2169 6506 2203
rect 6564 2169 6598 2203
rect 3260 1957 3330 2067
rect 3719 1804 3783 1872
rect 80 1724 114 1758
rect 208 1724 242 1758
rect 336 1724 370 1758
rect 464 1724 498 1758
rect 592 1724 626 1758
rect 720 1724 754 1758
rect 848 1724 882 1758
rect 976 1724 1010 1758
rect 1104 1724 1138 1758
rect 1232 1724 1266 1758
rect 1360 1724 1394 1758
rect 1488 1724 1522 1758
rect 1616 1724 1650 1758
rect 1744 1724 1778 1758
rect 1872 1724 1906 1758
rect 2000 1724 2034 1758
rect 2128 1724 2162 1758
rect 2256 1724 2290 1758
rect 2384 1724 2418 1758
rect 2512 1724 2546 1758
rect 2640 1724 2674 1758
rect 2768 1724 2802 1758
rect 2896 1724 2930 1758
rect 3024 1724 3058 1758
rect 3152 1724 3186 1758
rect 3280 1724 3314 1758
rect 3408 1724 3442 1758
rect 3536 1724 3570 1758
rect 3664 1724 3698 1758
rect 3792 1724 3826 1758
rect 3920 1724 3954 1758
rect 4048 1724 4082 1758
rect 4176 1724 4210 1758
rect 4304 1724 4338 1758
rect 4432 1724 4466 1758
rect 4560 1724 4594 1758
rect 4688 1724 4722 1758
rect 4816 1724 4850 1758
rect 4944 1724 4978 1758
rect 5072 1724 5106 1758
rect 5200 1724 5234 1758
rect 5328 1724 5362 1758
rect 5456 1724 5490 1758
rect 5584 1724 5618 1758
rect 5712 1724 5746 1758
rect 5840 1724 5874 1758
rect 5968 1724 6002 1758
rect 6096 1724 6130 1758
rect 6289 1625 6323 1659
rect 81 1526 115 1560
rect 209 1526 243 1560
rect 337 1526 371 1560
rect 465 1526 499 1560
rect 593 1526 627 1560
rect 721 1526 755 1560
rect 849 1526 883 1560
rect 977 1526 1011 1560
rect 1105 1526 1139 1560
rect 1233 1526 1267 1560
rect 1361 1526 1395 1560
rect 1489 1526 1523 1560
rect 1617 1526 1651 1560
rect 1745 1526 1779 1560
rect 1873 1526 1907 1560
rect 2001 1526 2035 1560
rect 2129 1526 2163 1560
rect 2257 1526 2291 1560
rect 2385 1526 2419 1560
rect 2513 1526 2547 1560
rect 2641 1526 2675 1560
rect 2769 1526 2803 1560
rect 2897 1526 2931 1560
rect 3025 1526 3059 1560
rect 3260 1424 3330 1480
rect 3875 1452 3909 1486
rect 4003 1452 4037 1486
rect 4131 1452 4165 1486
rect 4259 1452 4293 1486
rect 4387 1452 4421 1486
rect 4515 1452 4549 1486
rect 4643 1452 4677 1486
rect 4771 1452 4805 1486
rect 4899 1452 4933 1486
rect 5027 1452 5061 1486
rect 5155 1452 5189 1486
rect 5283 1452 5317 1486
rect 5535 1306 5569 1340
rect 5663 1306 5697 1340
rect 5791 1306 5825 1340
rect 5919 1306 5953 1340
rect 6047 1306 6081 1340
rect 6175 1306 6209 1340
rect 76 871 242 923
rect 3260 766 3330 833
rect 6565 537 6599 571
rect 3260 299 3330 366
rect 76 209 242 261
<< metal1 >>
rect 4 2203 6628 2234
rect 4 2169 33 2203
rect 67 2169 125 2203
rect 159 2169 217 2203
rect 251 2169 309 2203
rect 343 2169 401 2203
rect 435 2169 493 2203
rect 527 2169 585 2203
rect 619 2169 677 2203
rect 711 2169 769 2203
rect 803 2169 861 2203
rect 895 2169 953 2203
rect 987 2169 1045 2203
rect 1079 2169 1137 2203
rect 1171 2169 1229 2203
rect 1263 2169 1321 2203
rect 1355 2169 1413 2203
rect 1447 2169 1504 2203
rect 1538 2169 1596 2203
rect 1630 2169 1688 2203
rect 1722 2169 1780 2203
rect 1814 2169 1872 2203
rect 1906 2169 1964 2203
rect 1998 2169 2056 2203
rect 2090 2169 2148 2203
rect 2182 2169 2240 2203
rect 2274 2169 2332 2203
rect 2366 2169 2424 2203
rect 2458 2169 2516 2203
rect 2550 2169 2608 2203
rect 2642 2169 2700 2203
rect 2734 2169 2792 2203
rect 2826 2169 2884 2203
rect 2918 2169 2976 2203
rect 3010 2169 3068 2203
rect 3102 2169 3160 2203
rect 3194 2169 3252 2203
rect 3286 2169 3344 2203
rect 3378 2169 3436 2203
rect 3470 2169 3528 2203
rect 3562 2169 3620 2203
rect 3654 2169 3712 2203
rect 3746 2169 3804 2203
rect 3838 2169 3896 2203
rect 3930 2169 3988 2203
rect 4022 2169 4080 2203
rect 4114 2169 4172 2203
rect 4206 2169 4264 2203
rect 4298 2169 4356 2203
rect 4390 2169 4448 2203
rect 4482 2169 4540 2203
rect 4574 2169 4632 2203
rect 4666 2169 4724 2203
rect 4758 2169 4816 2203
rect 4850 2169 4908 2203
rect 4942 2169 5000 2203
rect 5034 2169 5092 2203
rect 5126 2169 5184 2203
rect 5218 2169 5276 2203
rect 5310 2169 5368 2203
rect 5402 2169 5460 2203
rect 5494 2169 5552 2203
rect 5586 2169 5644 2203
rect 5678 2169 5736 2203
rect 5770 2169 5828 2203
rect 5862 2169 5920 2203
rect 5954 2169 6012 2203
rect 6046 2169 6104 2203
rect 6138 2169 6196 2203
rect 6230 2169 6288 2203
rect 6322 2169 6380 2203
rect 6414 2169 6472 2203
rect 6506 2169 6564 2203
rect 6598 2169 6628 2203
rect 4 2138 6628 2169
rect 3254 2067 3336 2079
rect 3250 1957 3260 2067
rect 3330 1957 3340 2067
rect 3254 1945 3336 1957
rect 3713 1872 3789 1884
rect 3709 1801 3719 1872
rect 3783 1801 3793 1872
rect 3713 1792 3789 1801
rect 4 1758 6628 1764
rect 4 1724 80 1758
rect 114 1724 208 1758
rect 242 1724 336 1758
rect 370 1724 464 1758
rect 498 1724 592 1758
rect 626 1724 720 1758
rect 754 1724 848 1758
rect 882 1724 976 1758
rect 1010 1724 1104 1758
rect 1138 1724 1232 1758
rect 1266 1724 1360 1758
rect 1394 1724 1488 1758
rect 1522 1724 1616 1758
rect 1650 1724 1744 1758
rect 1778 1724 1872 1758
rect 1906 1724 2000 1758
rect 2034 1724 2128 1758
rect 2162 1724 2256 1758
rect 2290 1724 2384 1758
rect 2418 1724 2512 1758
rect 2546 1724 2640 1758
rect 2674 1724 2768 1758
rect 2802 1724 2896 1758
rect 2930 1724 3024 1758
rect 3058 1724 3152 1758
rect 3186 1724 3280 1758
rect 3314 1724 3408 1758
rect 3442 1724 3536 1758
rect 3570 1724 3664 1758
rect 3698 1724 3792 1758
rect 3826 1724 3920 1758
rect 3954 1724 4048 1758
rect 4082 1724 4176 1758
rect 4210 1724 4304 1758
rect 4338 1724 4432 1758
rect 4466 1724 4560 1758
rect 4594 1724 4688 1758
rect 4722 1724 4816 1758
rect 4850 1724 4944 1758
rect 4978 1724 5072 1758
rect 5106 1724 5200 1758
rect 5234 1724 5328 1758
rect 5362 1724 5456 1758
rect 5490 1724 5584 1758
rect 5618 1724 5712 1758
rect 5746 1724 5840 1758
rect 5874 1724 5968 1758
rect 6002 1724 6096 1758
rect 6130 1724 6628 1758
rect 4 1718 6628 1724
rect 6260 1659 6352 1690
rect 6260 1625 6289 1659
rect 6323 1625 6352 1659
rect 6260 1594 6352 1625
rect 5 1560 6628 1566
rect 5 1526 81 1560
rect 115 1526 209 1560
rect 243 1526 337 1560
rect 371 1526 465 1560
rect 499 1526 593 1560
rect 627 1526 721 1560
rect 755 1526 849 1560
rect 883 1526 977 1560
rect 1011 1526 1105 1560
rect 1139 1526 1233 1560
rect 1267 1526 1361 1560
rect 1395 1526 1489 1560
rect 1523 1526 1617 1560
rect 1651 1526 1745 1560
rect 1779 1526 1873 1560
rect 1907 1526 2001 1560
rect 2035 1526 2129 1560
rect 2163 1526 2257 1560
rect 2291 1526 2385 1560
rect 2419 1526 2513 1560
rect 2547 1526 2641 1560
rect 2675 1526 2769 1560
rect 2803 1526 2897 1560
rect 2931 1526 3025 1560
rect 3059 1526 6628 1560
rect 5 1520 6628 1526
rect 5 1446 3226 1492
rect 5 1372 3152 1418
rect 3106 1310 3152 1372
rect 3180 1384 3226 1446
rect 3254 1480 3336 1492
rect 3254 1412 3260 1480
rect 3330 1412 3336 1480
rect 3364 1486 6628 1492
rect 3364 1452 3875 1486
rect 3909 1452 4003 1486
rect 4037 1452 4131 1486
rect 4165 1452 4259 1486
rect 4293 1452 4387 1486
rect 4421 1452 4515 1486
rect 4549 1452 4643 1486
rect 4677 1452 4771 1486
rect 4805 1452 4899 1486
rect 4933 1452 5027 1486
rect 5061 1452 5155 1486
rect 5189 1452 5283 1486
rect 5317 1452 6628 1486
rect 3364 1446 6628 1452
rect 3364 1384 3410 1446
rect 3180 1338 3410 1384
rect 6181 1372 6628 1418
rect 6181 1346 6227 1372
rect 3471 1340 6227 1346
rect 3471 1310 5535 1340
rect 3106 1306 5535 1310
rect 5569 1306 5663 1340
rect 5697 1306 5791 1340
rect 5825 1306 5919 1340
rect 5953 1306 6047 1340
rect 6081 1306 6175 1340
rect 6209 1306 6227 1340
rect 3106 1300 6227 1306
rect 3106 1264 3517 1300
rect 3700 1249 6628 1270
rect 3700 1230 3719 1249
rect 3256 1174 3266 1230
rect 3330 1174 3340 1230
rect 3709 1193 3719 1230
rect 3783 1193 6628 1249
rect 3752 1174 6628 1193
rect 2 923 254 929
rect 2 871 76 923
rect 242 871 254 923
rect 2 865 254 871
rect 3248 833 3342 839
rect 3248 766 3260 833
rect 3330 766 3342 833
rect 3248 760 3342 766
rect 6536 571 6628 602
rect 6536 537 6565 571
rect 6599 537 6628 571
rect 6536 506 6628 537
rect 3248 366 3342 372
rect 3248 299 3260 366
rect 3330 299 3342 366
rect 3248 293 3342 299
rect 64 261 254 267
rect 64 209 76 261
rect 242 209 254 261
rect 64 203 254 209
<< via1 >>
rect 3260 1957 3330 2067
rect 3719 1804 3783 1872
rect 3719 1801 3783 1804
rect 3260 1424 3330 1480
rect 3260 1412 3330 1424
rect 3266 1174 3330 1230
rect 3719 1193 3783 1249
rect 76 871 242 923
rect 3260 766 3330 833
rect 3260 299 3330 366
rect 76 209 242 261
<< metal2 >>
rect 3260 2067 3330 2073
rect 3260 1480 3330 1957
rect 3260 1230 3330 1412
rect 3260 1174 3266 1230
rect 3719 1872 3783 1882
rect 3719 1249 3783 1801
rect 3719 1183 3783 1193
rect 76 923 242 933
rect 76 261 242 871
rect 3260 833 3330 1174
rect 3260 366 3330 766
rect 3260 289 3330 299
rect 76 199 242 209
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_0 ~/proj/pdk-installs-nbu/open-pdks-src/sky130/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1633901636
transform 1 0 4 0 1 10
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_1
timestamp 1633901636
transform 1 0 740 0 1 10
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_2
timestamp 1633901636
transform 1 0 1476 0 1 10
box -38 -48 774 592
use p-leg_fet_16  p-leg_fet_16_0
timestamp 1643073387
transform 1 0 1055 0 1 363
box -1089 -161 1089 198
use p-leg_fet_16  p-leg_fet_16_3
timestamp 1643073387
transform 1 0 1055 0 -1 769
box -1089 -161 1089 198
use p-leg_fet_16  p-leg_fet_16_1
timestamp 1643073387
transform 1 0 3103 0 1 363
box -1089 -161 1089 198
use p-leg_fet_16  p-leg_fet_16_4
timestamp 1643073387
transform 1 0 3103 0 -1 769
box -1089 -161 1089 198
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_3
timestamp 1633901636
transform 1 0 2212 0 1 10
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_4
timestamp 1633901636
transform 1 0 2948 0 1 10
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_5
timestamp 1633901636
transform 1 0 3684 0 1 10
box -38 -48 774 592
use p-leg_fet_16  p-leg_fet_16_2
timestamp 1643073387
transform 1 0 5151 0 1 363
box -1089 -161 1089 198
use p-leg_fet_16  p-leg_fet_16_5
timestamp 1643073387
transform 1 0 5151 0 -1 769
box -1089 -161 1089 198
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_6
timestamp 1633901636
transform 1 0 4420 0 1 10
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_7
timestamp 1633901636
transform 1 0 5156 0 1 10
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_8
timestamp 1633901636
transform 1 0 5892 0 1 10
box -38 -48 774 592
use p-leg_6  p-leg_6_2
timestamp 1643158822
transform 1 0 2594 0 -1 1415
box -1089 -161 -191 198
use p-leg_6  p-leg_6_1
timestamp 1643158822
transform 1 0 1826 0 -1 1415
box -1089 -161 -191 198
use p-leg_6  p-leg_6_0
timestamp 1643158822
transform 1 0 1058 0 -1 1415
box -1089 -161 -191 198
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_10
timestamp 1633901636
transform 1 0 740 0 1 1098
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_9
timestamp 1633901636
transform 1 0 4 0 1 1098
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_11
timestamp 1633901636
transform 1 0 1476 0 1 1098
box -38 -48 774 592
use p-leg_6  p-leg_6_4
timestamp 1643158822
transform 1 0 4852 0 -1 1341
box -1089 -161 -191 198
use p-leg_6  p-leg_6_3
timestamp 1643158822
transform 1 0 3362 0 -1 1415
box -1089 -161 -191 198
use p-leg_polyres  p-leg_polyres_0
timestamp 1643152784
transform 0 -1 3515 1 0 1197
box -33 -253 33 253
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_13
timestamp 1633901636
transform 1 0 2948 0 1 1098
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_12
timestamp 1633901636
transform 1 0 2212 0 1 1098
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_14
timestamp 1633901636
transform 1 0 3684 0 1 1098
box -38 -48 774 592
use p-leg_6  p-leg_6_5
timestamp 1643158822
transform 1 0 5620 0 -1 1341
box -1089 -161 -191 198
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_16
timestamp 1633901636
transform 1 0 5156 0 1 1098
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_15
timestamp 1633901636
transform 1 0 4420 0 1 1098
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  sky130_fd_sc_hd__fill_8_17
timestamp 1633901636
transform 1 0 5892 0 1 1098
box -38 -48 774 592
use p-leg_fet_16  p-leg_fet_16_6
timestamp 1643073387
transform -1 0 3105 0 1 1869
box -1089 -161 1089 198
use p-leg_fet_16  p-leg_fet_16_8
timestamp 1643073387
transform -1 0 1057 0 1 1869
box -1089 -161 1089 198
use p-leg_fet_16  p-leg_fet_16_7
timestamp 1643073387
transform -1 0 5153 0 1 1869
box -1089 -161 1089 198
use p-leg_6  p-leg_6_6
timestamp 1643158822
transform 1 0 6512 0 1 1451
box -1089 -161 -191 198
<< labels >>
flabel metal1 s 40 895 40 895 7 FreeSerif 640 0 0 0 n_pu_ctrl
port 1 w
flabel metal1 s 6586 1220 6586 1220 3 FreeSerif 640 0 0 0 DQ
port 2 e
flabel metal1 s 30 553 30 553 7 FreeSerif 640 0 0 0 VDD
port 3 w
flabel metal1 s 30 1641 30 1641 7 FreeSerif 640 0 0 0 VDD
port 3 w
flabel metal1 s 26 1740 26 1740 7 FreeSerif 640 0 0 0 n_cal_ctrl[0]
port 4 w
flabel metal1 s 27 1542 27 1542 7 FreeSerif 640 0 0 0 n_cal_ctrl[1]
port 5 w
flabel metal1 s 27 1468 27 1468 7 FreeSerif 640 0 0 0 n_cal_ctrl[2]
port 6 w
flabel metal1 s 27 1394 27 1394 7 FreeSerif 640 0 0 0 n_cal_ctrl[3]
port 7 w
flabel metal1 3294 997 3294 997 7 FreeSerif 640 0 0 0 v_pullup
<< end >>
