* Fast-Fast corner (ff)
.lib ff
.param mc_mm_switch=0
.param mc_pr_switch=0
* MOSFET
.include "sky130_libs/corners/ff.spice"
* Resistor/Capacitor
.include "sky130_libs/r+c/res_typical__cap_typical.spice"
.include "sky130_libs/r+c/res_typical__cap_typical__lin.spice"
* Special cells
.include "sky130_libs/corners/ff/specialized_cells.spice"
.endl ff
