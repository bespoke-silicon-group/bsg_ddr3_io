**.subckt p-leg_tb
Vctrl0 VDD n_cal_ctrl[0] SED_vctrl0_SED
Vctrl1 VDD n_cal_ctrl[1] SED_vctrl1_SED
Vctrl2 VDD n_cal_ctrl[2] SED_vctrl2_SED
Vctrl3 VDD n_cal_ctrl[3] SED_vctrl3_SED
Vgate VDD n_pu_ctrl SED_vg_SED
Vtest DQ VDDQ 0
.save  i(vtest)
Vpinvoltage v1v5 VDDQ 0
X1 DQ n_pu_ctrl n_cal_ctrl[3] n_cal_ctrl[2] n_cal_ctrl[1] n_cal_ctrl[0] p-leg
**** begin user architecture code
 ** Local library links to pdk
.lib ./sky130/libs/SED_process_SED_lib.spice SED_process_SED

**** end user architecture code
**.ends

* expanding   symbol:  p-leg.sym # of pins=3
* sym_path: /mnt/users/ssd2/homes/hinesd3/proj/sstl-design/schem/p-leg.sym
* sch_path: /mnt/users/ssd2/homes/hinesd3/proj/sstl-design/schem/p-leg.sch
.subckt p-leg  DQ  n_pu_ctrl  n_cal_ctrl[3] n_cal_ctrl[2] n_cal_ctrl[1] n_cal_ctrl[0]
*.ipin n_cal_ctrl[3],n_cal_ctrl[2],n_cal_ctrl[1],n_cal_ctrl[0]
*.ipin n_pu_ctrl
*.iopin DQ
R1 DQ net1 sky130_fd_pr__res_generic_po W=0.33 L=1.8 m=1
XMpullup net1 n_pu_ctrl VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=96 m=96
XMctrl0 DQ n_cal_ctrl[0] net1 VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=48 m=48
XMctrl1 DQ n_cal_ctrl[1] net1 VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=24 m=24
XMctrl2 DQ n_cal_ctrl[2] net1 VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=12 m=12
XMctrl3 DQ n_cal_ctrl[3] net1 VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=6 m=6
.ends

.GLOBAL VDD
**** begin user architecture code



* power voltage
vvdd VDD 0 SED_vdd_SED
vv1v5 v1v5 0 1.5

.control
save all
set temp=SED_temp_SED

* RUN SIMULATION
dc Vpinvoltage 0.3 1.2 0.05
* OUTPUT
print (SED_vdd_SED-vddq)/i(vtest)
wrdata out/SED_plotName_SED/SED_plotName_SED.txt (SED_vdd_SED-vddq)/i(vtest)
set hcopydevtype = svg
hardcopy ./out/SED_plotName_SED/SED_plotName_SED.svg (SED_vdd_SED-vddq)/I(vtest) vs vddq title 'Resistance vs pin voltage'

.endc


**** end user architecture code
.end
