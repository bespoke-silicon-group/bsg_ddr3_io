* High-Low corner with mismatch (hl_mm)
.lib hl_mm
.param mc_mm_switch=1
.param mc_pr_switch=0
* MOSFET
.include "sky130_libs/corners/tt.spice"
* Resistor/Capacitor
.include "sky130_libs/r+c/res_high__cap_low.spice"
.include "sky130_libs/r+c/res_high__cap_low__lin.spice"
* Special cells
.include "sky130_libs/corners/tt/specialized_cells.spice"
.endl hl_mm
