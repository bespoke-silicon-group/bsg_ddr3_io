* Fast-Fast corner with mismatch (ff_mm)
.lib ff_mm
.param mc_mm_switch=1
.param mc_pr_switch=0
* MOSFET
.include "sky130_libs/corners/ff.spice"
* Resistor/Capacitor
.include "sky130_libs/r+c/res_typical__cap_typical.spice"
.include "sky130_libs/r+c/res_typical__cap_typical__lin.spice"
* Special cells
.include "sky130_libs/corners/ff/specialized_cells.spice"
.endl ff_mm
