magic
tech sky130A
magscale 1 2
timestamp 1643073387
<< nwell >>
rect -1089 -100 1089 198
<< pmoslvt >>
rect -995 -64 -925 136
rect -867 -64 -797 136
rect -739 -64 -669 136
rect -611 -64 -541 136
rect -483 -64 -413 136
rect -355 -64 -285 136
rect -227 -64 -157 136
rect -99 -64 -29 136
rect 29 -64 99 136
rect 157 -64 227 136
rect 285 -64 355 136
rect 413 -64 483 136
rect 541 -64 611 136
rect 669 -64 739 136
rect 797 -64 867 136
rect 925 -64 995 136
<< pdiff >>
rect -1053 124 -995 136
rect -1053 53 -1041 124
rect -1007 53 -995 124
rect -1053 -64 -995 53
rect -925 19 -867 136
rect -925 -52 -913 19
rect -879 -52 -867 19
rect -925 -64 -867 -52
rect -797 124 -739 136
rect -797 53 -785 124
rect -751 53 -739 124
rect -797 -64 -739 53
rect -669 19 -611 136
rect -669 -52 -657 19
rect -623 -52 -611 19
rect -669 -64 -611 -52
rect -541 124 -483 136
rect -541 53 -529 124
rect -495 53 -483 124
rect -541 -64 -483 53
rect -413 19 -355 136
rect -413 -52 -401 19
rect -367 -52 -355 19
rect -413 -64 -355 -52
rect -285 124 -227 136
rect -285 53 -273 124
rect -239 53 -227 124
rect -285 -64 -227 53
rect -157 19 -99 136
rect -157 -52 -145 19
rect -111 -52 -99 19
rect -157 -64 -99 -52
rect -29 124 29 136
rect -29 53 -17 124
rect 17 53 29 124
rect -29 -64 29 53
rect 99 19 157 136
rect 99 -52 111 19
rect 145 -52 157 19
rect 99 -64 157 -52
rect 227 124 285 136
rect 227 53 239 124
rect 273 53 285 124
rect 227 -64 285 53
rect 355 19 413 136
rect 355 -52 367 19
rect 401 -52 413 19
rect 355 -64 413 -52
rect 483 124 541 136
rect 483 53 495 124
rect 529 53 541 124
rect 483 -64 541 53
rect 611 19 669 136
rect 611 -52 623 19
rect 657 -52 669 19
rect 611 -64 669 -52
rect 739 124 797 136
rect 739 53 751 124
rect 785 53 797 124
rect 739 -64 797 53
rect 867 19 925 136
rect 867 -52 879 19
rect 913 -52 925 19
rect 867 -64 925 -52
rect 995 124 1053 136
rect 995 53 1007 124
rect 1041 53 1053 124
rect 995 -64 1053 53
<< pdiffc >>
rect -1041 53 -1007 124
rect -913 -52 -879 19
rect -785 53 -751 124
rect -657 -52 -623 19
rect -529 53 -495 124
rect -401 -52 -367 19
rect -273 53 -239 124
rect -145 -52 -111 19
rect -17 53 17 124
rect 111 -52 145 19
rect 239 53 273 124
rect 367 -52 401 19
rect 495 53 529 124
rect 623 -52 657 19
rect 751 53 785 124
rect 879 -52 913 19
rect 1007 53 1041 124
<< poly >>
rect -995 136 -925 162
rect -867 136 -797 162
rect -739 136 -669 162
rect -611 136 -541 162
rect -483 136 -413 162
rect -355 136 -285 162
rect -227 136 -157 162
rect -99 136 -29 162
rect 29 136 99 162
rect 157 136 227 162
rect 285 136 355 162
rect 413 136 483 162
rect 541 136 611 162
rect 669 136 739 162
rect 797 136 867 162
rect 925 136 995 162
rect -995 -79 -925 -64
rect -867 -79 -797 -64
rect -739 -79 -669 -64
rect -611 -79 -541 -64
rect -483 -79 -413 -64
rect -355 -79 -285 -64
rect -227 -79 -157 -64
rect -99 -79 -29 -64
rect 29 -79 99 -64
rect 157 -79 227 -64
rect 285 -79 355 -64
rect 413 -79 483 -64
rect 541 -79 611 -64
rect 669 -79 739 -64
rect 797 -79 867 -64
rect 925 -79 995 -64
rect -1053 -111 1053 -79
rect -1053 -145 -979 -111
rect -941 -145 -851 -111
rect -813 -145 -723 -111
rect -685 -145 -595 -111
rect -557 -145 -467 -111
rect -429 -145 -339 -111
rect -301 -145 -211 -111
rect -173 -145 -83 -111
rect -45 -145 45 -111
rect 83 -145 173 -111
rect 211 -145 301 -111
rect 339 -145 429 -111
rect 467 -145 557 -111
rect 595 -145 685 -111
rect 723 -145 813 -111
rect 851 -145 941 -111
rect 979 -145 1053 -111
rect -1053 -161 1053 -145
<< polycont >>
rect -979 -145 -941 -111
rect -851 -145 -813 -111
rect -723 -145 -685 -111
rect -595 -145 -557 -111
rect -467 -145 -429 -111
rect -339 -145 -301 -111
rect -211 -145 -173 -111
rect -83 -145 -45 -111
rect 45 -145 83 -111
rect 173 -145 211 -111
rect 301 -145 339 -111
rect 429 -145 467 -111
rect 557 -145 595 -111
rect 685 -145 723 -111
rect 813 -145 851 -111
rect 941 -145 979 -111
<< locali >>
rect -1041 124 -1007 198
rect -1041 37 -1007 53
rect -785 124 -751 198
rect -913 19 -879 52
rect -785 37 -751 53
rect -529 124 -495 198
rect -1041 -52 -913 3
rect -657 19 -623 52
rect -529 37 -495 53
rect -273 124 -239 198
rect -879 -52 -657 3
rect -401 19 -367 52
rect -273 37 -239 53
rect -17 124 17 198
rect -623 -52 -401 3
rect -145 19 -111 52
rect -17 37 17 53
rect 239 124 273 198
rect -367 -52 -145 3
rect 111 19 145 52
rect 239 37 273 53
rect 495 124 529 198
rect -111 -52 111 3
rect 367 19 401 52
rect 495 37 529 53
rect 751 124 785 198
rect 145 -52 367 3
rect 623 19 657 52
rect 751 37 785 53
rect 1007 124 1041 198
rect 401 -52 623 3
rect 879 19 913 52
rect 1007 37 1041 53
rect 657 -52 879 3
rect 913 -52 1041 3
rect -1041 -68 1041 -52
rect -1053 -145 -979 -111
rect -941 -145 -851 -111
rect -813 -145 -723 -111
rect -685 -145 -595 -111
rect -557 -145 -467 -111
rect -429 -145 -339 -111
rect -301 -145 -211 -111
rect -173 -145 -83 -111
rect -45 -145 45 -111
rect 83 -145 173 -111
rect 211 -145 301 -111
rect 339 -145 429 -111
rect 467 -145 557 -111
rect 595 -145 685 -111
rect 723 -145 813 -111
rect 851 -145 941 -111
rect 979 -145 1053 -111
<< properties >>
string gencell sky130_fd_pr__pfet_01v8_lvt
string parameters w 1.0 l 0.35 m 1 nf 16 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
string library sky130
<< end >>
